module RiscvTrans(
  input  [31:0] io_inst, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input         io_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output        io_mem_read_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_mem_read_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [6:0]  io_mem_read_memWidth, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_mem_read_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output        io_mem_write_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_mem_write_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [6:0]  io_mem_write_memWidth, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_mem_write_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_4, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_5, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_6, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_7, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_8, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_9, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_10, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_11, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_12, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_13, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_14, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_15, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_16, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_17, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_18, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_19, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_20, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_21, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_22, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_23, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_24, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_25, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_26, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_27, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_28, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_29, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_30, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_31, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_pc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_misa, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mvendorid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_marchid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mimpid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mhartid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mstatus, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mtvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mcounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_medeleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mip, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mie, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mcause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mtval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_scause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_stvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_sepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [7:0]  io_now_csr_MXLEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [1:0]  io_now_internal_privilegeMode, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_4, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_5, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_6, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_7, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_8, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_9, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_10, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_11, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_12, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_13, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_14, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_15, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_16, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_17, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_18, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_19, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_20, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_21, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_22, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_23, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_24, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_25, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_26, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_27, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_28, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_29, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_30, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_31, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_pc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_misa, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mvendorid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_marchid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mimpid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mhartid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mstatus, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mtvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mcounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_medeleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mip, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mie, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mcause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mtval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_scause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_stvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_sepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [7:0]  io_next_csr_MXLEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [1:0]  io_next_internal_privilegeMode, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output        io_event_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_event_cause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_event_exceptionPC, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_event_exceptionInst // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
);
  wire [31:0] inst = io_valid ? io_inst : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 130:16 112:21]
  wire [31:0] _T_656 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_657 = 32'h3003 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _T_1144 = inst & 32'hfe007fff; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1145 = 32'h12000073 == _T_1144; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1139 = 32'h10500073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1132 = 32'h30200073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1125 = 32'h10200073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _T_1117 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1118 = 32'h200703b == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1111 = 32'h200603b == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1104 = 32'h200503b == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1097 = 32'h200403b == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1090 = 32'h200003b == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1083 = 32'h2007033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1076 = 32'h2006033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1069 = 32'h2005033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1062 = 32'h2004033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1055 = 32'h2003033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1048 = 32'h2002033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1041 = 32'h2001033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1034 = 32'h2000033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _T_1007 = inst & 32'he003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_1010 = inst[11:7] != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:63]
  wire  _T_1011 = 32'h2001 == _T_1007 & _T_1010; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_971 = 32'h6002 == _T_1007 & _T_1010; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [31:0] _T_960 = inst & 32'hef83; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_961 = 32'h1 == _T_960; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _T_916 = inst & 32'hf003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_922 = _T_1010 & inst[6:2] != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 76:105]
  wire  _T_923 = 32'h9002 == _T_916 & _T_922; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_911 = 32'h8002 == _T_916 & _T_922; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [5:0] _T_858 = {inst[12],inst[6:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:14]
  wire  _T_859 = _T_858 != 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:37]
  wire  _T_861 = _T_1010 & _T_859; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 65:105]
  wire  _T_862 = 32'h2 == _T_1007 & _T_861; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_836 = 32'h6101 == _T_960 & _T_859; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_824 = 32'h1 == _T_1007 & _T_861; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_808 = _T_1010 & inst[11:7] != 5'h2 & _T_859; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 44:130]
  wire  _T_809 = 32'h6001 == _T_1007 & _T_808; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_791 = 32'h4001 == _T_1007 & _T_1010; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [31:0] _T_760 = inst & 32'hf07f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_764 = 32'h9002 == _T_760 & _T_1010; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_755 = 32'h8002 == _T_760 & _T_1010; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_704 = 32'h4002 == _T_1007 & _T_1010; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_677 = 32'h3023 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_637 = 32'h6003 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_630 = 32'h4000503b == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_623 = 32'h4000003b == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_616 = 32'h503b == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_609 = 32'h103b == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_602 = 32'h3b == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_595 = 32'h40005033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_588 = 32'h5033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_581 = 32'h1033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_575 = 32'h4000501b == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_569 = 32'h501b == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_563 = 32'h101b == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _T_556 = inst & 32'hfc00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_557 = 32'h40005013 == _T_556; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_551 = 32'h5013 == _T_556; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_545 = 32'h1013 == _T_556; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_539 = 32'h1b == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_533 = 32'hf == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_524 = 32'h73 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_518 = 32'h100073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_494 = 32'h2023 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_470 = 32'h1023 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_447 = 32'h23 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_427 = 32'h5003 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_408 = 32'h4003 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_388 = 32'h2003 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_368 = 32'h1003 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_348 = 32'h3 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_321 = 32'h7063 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_292 = 32'h5063 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_265 = 32'h6063 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_236 = 32'h4063 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_209 = 32'h1063 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_182 = 32'h63 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_157 = 32'h67 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_119 = 32'h40000033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_98 = 32'h4033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_91 = 32'h6033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_84 = 32'h7033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_77 = 32'h3033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_70 = 32'h2033 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_63 = 32'h33 == _T_1117; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_31 = 32'h4013 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_25 = 32'h6013 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_19 = 32'h7013 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_13 = 32'h3013 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_7 = 32'h2013 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1 = 32'h13 == _T_656; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [4:0] _GEN_66 = _T_1 ? inst[19:15] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 19:24]
  wire [4:0] _GEN_137 = _T_7 ? inst[19:15] : _GEN_66; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_208 = _T_13 ? inst[19:15] : _GEN_137; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_279 = _T_19 ? inst[19:15] : _GEN_208; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_350 = _T_25 ? inst[19:15] : _GEN_279; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_421 = _T_31 ? inst[19:15] : _GEN_350; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_492 = _T_545 ? inst[19:15] : _GEN_421; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_563 = _T_551 ? inst[19:15] : _GEN_492; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_634 = _T_557 ? inst[19:15] : _GEN_563; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_876 = _T_63 ? inst[19:15] : _GEN_634; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_947 = _T_70 ? inst[19:15] : _GEN_876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1018 = _T_77 ? inst[19:15] : _GEN_947; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1089 = _T_84 ? inst[19:15] : _GEN_1018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1160 = _T_91 ? inst[19:15] : _GEN_1089; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1231 = _T_98 ? inst[19:15] : _GEN_1160; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1302 = _T_581 ? inst[19:15] : _GEN_1231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1373 = _T_588 ? inst[19:15] : _GEN_1302; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1444 = _T_119 ? inst[19:15] : _GEN_1373; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1515 = _T_595 ? inst[19:15] : _GEN_1444; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1736 = _T_157 ? inst[19:15] : _GEN_1515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1792 = _T_182 ? inst[19:15] : _GEN_1736; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1817 = _T_209 ? inst[19:15] : _GEN_1792; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1842 = _T_236 ? inst[19:15] : _GEN_1817; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1867 = _T_265 ? inst[19:15] : _GEN_1842; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1892 = _T_292 ? inst[19:15] : _GEN_1867; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1917 = _T_321 ? inst[19:15] : _GEN_1892; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1999 = _T_348 ? inst[19:15] : _GEN_1917; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2112 = _T_368 ? inst[19:15] : _GEN_1999; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2225 = _T_388 ? inst[19:15] : _GEN_2112; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2303 = _T_408 ? inst[19:15] : _GEN_2225; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2416 = _T_427 ? inst[19:15] : _GEN_2303; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2463 = _T_447 ? inst[19:15] : _GEN_2416; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2483 = _T_470 ? inst[19:15] : _GEN_2463; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2503 = _T_494 ? inst[19:15] : _GEN_2483; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2516 = _T_518 ? inst[19:15] : _GEN_2503; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2534 = _T_524 ? inst[19:15] : _GEN_2516; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2545 = _T_533 ? inst[19:15] : _GEN_2534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2584 = _T_539 ? inst[19:15] : _GEN_2545; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2655 = _T_545 ? inst[19:15] : _GEN_2584; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2726 = _T_551 ? inst[19:15] : _GEN_2655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2797 = _T_557 ? inst[19:15] : _GEN_2726; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2868 = _T_563 ? inst[19:15] : _GEN_2797; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2939 = _T_569 ? inst[19:15] : _GEN_2868; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3010 = _T_575 ? inst[19:15] : _GEN_2939; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3082 = _T_581 ? inst[19:15] : _GEN_3010; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3153 = _T_588 ? inst[19:15] : _GEN_3082; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3224 = _T_595 ? inst[19:15] : _GEN_3153; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3295 = _T_602 ? inst[19:15] : _GEN_3224; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3366 = _T_609 ? inst[19:15] : _GEN_3295; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3437 = _T_616 ? inst[19:15] : _GEN_3366; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3508 = _T_623 ? inst[19:15] : _GEN_3437; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3579 = _T_630 ? inst[19:15] : _GEN_3508; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3686 = _T_637 ? inst[19:15] : _GEN_3579; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3799 = _T_657 ? inst[19:15] : _GEN_3686; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3850 = _T_677 ? inst[19:15] : _GEN_3799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3896 = _T_704 ? inst[11:7] : _GEN_3850; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4146 = _T_755 ? inst[11:7] : _GEN_3896; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4154 = _T_764 ? inst[11:7] : _GEN_4146; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4284 = _T_791 ? inst[11:7] : _GEN_4154; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4356 = _T_809 ? inst[11:7] : _GEN_4284; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4459 = _T_824 ? inst[11:7] : _GEN_4356; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4498 = _T_836 ? inst[11:7] : _GEN_4459; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 220:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4607 = _T_862 ? inst[11:7] : _GEN_4498; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4990 = _T_911 ? inst[11:7] : _GEN_4607; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5060 = _T_923 ? inst[11:7] : _GEN_4990; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5639 = _T_961 ? inst[11:7] : _GEN_5060; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 259:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5678 = _T_971 ? inst[11:7] : _GEN_5639; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5946 = _T_1011 ? inst[11:7] : _GEN_5678; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6288 = _T_1034 ? inst[19:15] : _GEN_5946; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6359 = _T_1041 ? inst[19:15] : _GEN_6288; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6430 = _T_1048 ? inst[19:15] : _GEN_6359; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6501 = _T_1055 ? inst[19:15] : _GEN_6430; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6572 = _T_1062 ? inst[19:15] : _GEN_6501; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6643 = _T_1069 ? inst[19:15] : _GEN_6572; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6714 = _T_1076 ? inst[19:15] : _GEN_6643; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6785 = _T_1083 ? inst[19:15] : _GEN_6714; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6856 = _T_1090 ? inst[19:15] : _GEN_6785; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6927 = _T_1097 ? inst[19:15] : _GEN_6856; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6998 = _T_1104 ? inst[19:15] : _GEN_6927; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7069 = _T_1111 ? inst[19:15] : _GEN_6998; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7140 = _T_1118 ? inst[19:15] : _GEN_7069; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7189 = _T_1125 ? inst[19:15] : _GEN_7140; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7210 = _T_1132 ? inst[19:15] : _GEN_7189; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7224 = _T_1139 ? inst[19:15] : _GEN_7210; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7231 = _T_1145 ? inst[19:15] : _GEN_7224; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] rs1 = io_valid ? _GEN_7231 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 19:24]
  wire [63:0] _GEN_1 = 5'h1 == rs1 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_2 = 5'h2 == rs1 ? io_now_reg_2 : _GEN_1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_3 = 5'h3 == rs1 ? io_now_reg_3 : _GEN_2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_4 = 5'h4 == rs1 ? io_now_reg_4 : _GEN_3; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_5 = 5'h5 == rs1 ? io_now_reg_5 : _GEN_4; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_6 = 5'h6 == rs1 ? io_now_reg_6 : _GEN_5; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_7 = 5'h7 == rs1 ? io_now_reg_7 : _GEN_6; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_8 = 5'h8 == rs1 ? io_now_reg_8 : _GEN_7; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_9 = 5'h9 == rs1 ? io_now_reg_9 : _GEN_8; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_10 = 5'ha == rs1 ? io_now_reg_10 : _GEN_9; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_11 = 5'hb == rs1 ? io_now_reg_11 : _GEN_10; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_12 = 5'hc == rs1 ? io_now_reg_12 : _GEN_11; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_13 = 5'hd == rs1 ? io_now_reg_13 : _GEN_12; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_14 = 5'he == rs1 ? io_now_reg_14 : _GEN_13; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_15 = 5'hf == rs1 ? io_now_reg_15 : _GEN_14; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_16 = 5'h10 == rs1 ? io_now_reg_16 : _GEN_15; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_17 = 5'h11 == rs1 ? io_now_reg_17 : _GEN_16; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_18 = 5'h12 == rs1 ? io_now_reg_18 : _GEN_17; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_19 = 5'h13 == rs1 ? io_now_reg_19 : _GEN_18; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_20 = 5'h14 == rs1 ? io_now_reg_20 : _GEN_19; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_21 = 5'h15 == rs1 ? io_now_reg_21 : _GEN_20; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_22 = 5'h16 == rs1 ? io_now_reg_22 : _GEN_21; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_23 = 5'h17 == rs1 ? io_now_reg_23 : _GEN_22; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_24 = 5'h18 == rs1 ? io_now_reg_24 : _GEN_23; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_25 = 5'h19 == rs1 ? io_now_reg_25 : _GEN_24; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_26 = 5'h1a == rs1 ? io_now_reg_26 : _GEN_25; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_27 = 5'h1b == rs1 ? io_now_reg_27 : _GEN_26; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_28 = 5'h1c == rs1 ? io_now_reg_28 : _GEN_27; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_29 = 5'h1d == rs1 ? io_now_reg_29 : _GEN_28; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_30 = 5'h1e == rs1 ? io_now_reg_30 : _GEN_29; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_31 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [11:0] _GEN_65 = _T_1 ? inst[31:20] : 12'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 38:27]
  wire [11:0] _GEN_136 = _T_7 ? inst[31:20] : _GEN_65; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_207 = _T_13 ? inst[31:20] : _GEN_136; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_278 = _T_19 ? inst[31:20] : _GEN_207; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_349 = _T_25 ? inst[31:20] : _GEN_278; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_420 = _T_31 ? inst[31:20] : _GEN_349; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_491 = _T_545 ? inst[31:20] : _GEN_420; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_562 = _T_551 ? inst[31:20] : _GEN_491; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_633 = _T_557 ? inst[31:20] : _GEN_562; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_1735 = _T_157 ? inst[31:20] : _GEN_633; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_1998 = _T_348 ? inst[31:20] : _GEN_1735; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2111 = _T_368 ? inst[31:20] : _GEN_1998; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2224 = _T_388 ? inst[31:20] : _GEN_2111; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2302 = _T_408 ? inst[31:20] : _GEN_2224; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2415 = _T_427 ? inst[31:20] : _GEN_2302; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2515 = _T_518 ? inst[31:20] : _GEN_2415; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2533 = _T_524 ? inst[31:20] : _GEN_2515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2544 = _T_533 ? inst[31:20] : _GEN_2533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2583 = _T_539 ? inst[31:20] : _GEN_2544; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2654 = _T_545 ? inst[31:20] : _GEN_2583; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2725 = _T_551 ? inst[31:20] : _GEN_2654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2796 = _T_557 ? inst[31:20] : _GEN_2725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2867 = _T_563 ? inst[31:20] : _GEN_2796; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2938 = _T_569 ? inst[31:20] : _GEN_2867; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_3009 = _T_575 ? inst[31:20] : _GEN_2938; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_3685 = _T_637 ? inst[31:20] : _GEN_3009; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_3798 = _T_657 ? inst[31:20] : _GEN_3685; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_7188 = _T_1125 ? inst[31:20] : _GEN_3798; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_7209 = _T_1132 ? inst[31:20] : _GEN_7188; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_7223 = _T_1139 ? inst[31:20] : _GEN_7209; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_7230 = _T_1145 ? inst[31:20] : _GEN_7223; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] imm_11_0 = io_valid ? _GEN_7230 : 12'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 38:27]
  wire  imm_signBit_50 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [51:0] _imm_T_320 = imm_signBit_50 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _imm_T_321 = {_imm_T_320,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [5:0] _imm_T_306 = {inst[12],inst[6],inst[5],inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  imm_signBit_46 = _imm_T_306[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [57:0] _imm_T_308 = imm_signBit_46 ? 58'h3ffffffffffffff : 58'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _imm_T_309 = {_imm_T_308,inst[12],inst[6],inst[5],inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  _T_996 = 32'he000 == _T_1007; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [63:0] _imm_T_299 = {56'h0,inst[6],inst[5],inst[12],inst[11],inst[10],3'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire  _T_987 = 32'h6000 == _T_1007; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_978 = 32'he002 == _T_1007; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [63:0] _imm_T_283 = {55'h0,inst[9],inst[8],inst[7],inst[12],inst[11],inst[10],3'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [63:0] _imm_T_274 = {55'h0,inst[4],inst[3],inst[2],inst[12],inst[6],inst[5],3'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _T_896 = inst & 32'hec03; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_897 = 32'h8801 == _T_896; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_889 = 32'h8401 == _T_896 & _T_859; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_875 = 32'h8001 == _T_896 & _T_859; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_779 = 32'he001 == _T_1007; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [8:0] _imm_T_221 = {inst[12],inst[6],inst[5],inst[2],inst[11],inst[10],inst[4],inst[3],1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire  imm_signBit_43 = _imm_T_221[8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [54:0] _imm_T_223 = imm_signBit_43 ? 55'h7fffffffffffff : 55'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _imm_T_224 = {_imm_T_223,inst[12],inst[6],inst[5],inst[2],inst[11],inst[10],inst[4],inst[3],1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  _T_770 = 32'hc001 == _T_1007; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [4:0] imm_lo_12 = {inst[2],inst[11],inst[5],inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [11:0] _imm_T_195 = {inst[12],inst[8],inst[10],inst[9],inst[6],inst[7],imm_lo_12,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire  imm_signBit_41 = _imm_T_195[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [51:0] _imm_T_197 = imm_signBit_41 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _imm_T_198 = {_imm_T_197,inst[12],inst[8],inst[10],inst[9],inst[6],inst[7],imm_lo_12,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  _T_741 = 32'ha001 == _T_1007; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_729 = 32'hc000 == _T_1007; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [63:0] _imm_T_166 = {57'h0,inst[5],inst[12],inst[11],inst[10],inst[6],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire  _T_720 = 32'h4000 == _T_1007; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_711 = 32'hc002 == _T_1007; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [63:0] _imm_T_150 = {56'h0,inst[8],inst[7],inst[12],inst[11],inst[10],inst[9],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [63:0] _imm_T_141 = {56'h0,inst[3],inst[2],inst[12],inst[6],inst[5],inst[4],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [6:0] _GEN_2461 = _T_447 ? inst[31:25] : 7'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:27]
  wire [6:0] _GEN_2481 = _T_470 ? inst[31:25] : _GEN_2461; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_2501 = _T_494 ? inst[31:25] : _GEN_2481; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_3848 = _T_677 ? inst[31:25] : _GEN_2501; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] imm_11_5 = io_valid ? _GEN_3848 : 7'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:27]
  wire [4:0] _GEN_2465 = _T_447 ? inst[11:7] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:62]
  wire [4:0] _GEN_2485 = _T_470 ? inst[11:7] : _GEN_2465; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2505 = _T_494 ? inst[11:7] : _GEN_2485; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3852 = _T_677 ? inst[11:7] : _GEN_2505; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] imm_4_0 = io_valid ? _GEN_3852 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:62]
  wire [11:0] _imm_T_129 = {imm_11_5,imm_4_0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:141]
  wire  imm_signBit_39 = _imm_T_129[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [51:0] _imm_T_131 = imm_signBit_39 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _imm_T_132 = {_imm_T_131,imm_11_5,imm_4_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  _GEN_1789 = _T_182 & inst[31]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:27]
  wire  _GEN_1814 = _T_209 ? inst[31] : _GEN_1789; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1839 = _T_236 ? inst[31] : _GEN_1814; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1864 = _T_265 ? inst[31] : _GEN_1839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1889 = _T_292 ? inst[31] : _GEN_1864; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1914 = _T_321 ? inst[31] : _GEN_1889; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  imm_12 = io_valid & _GEN_1914; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:27]
  wire [31:0] _T_132 = inst & 32'h7f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_133 = 32'h6f == _T_132; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _GEN_1623 = _T_133 & inst[20]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:132]
  wire  _GEN_1795 = _T_182 ? inst[7] : _GEN_1623; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1820 = _T_209 ? inst[7] : _GEN_1795; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1845 = _T_236 ? inst[7] : _GEN_1820; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1870 = _T_265 ? inst[7] : _GEN_1845; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1895 = _T_292 ? inst[7] : _GEN_1870; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1920 = _T_321 ? inst[7] : _GEN_1895; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  imm_11 = io_valid & _GEN_1920; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:132]
  wire [5:0] _GEN_1790 = _T_182 ? inst[30:25] : 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:62]
  wire [5:0] _GEN_1815 = _T_209 ? inst[30:25] : _GEN_1790; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_1840 = _T_236 ? inst[30:25] : _GEN_1815; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_1865 = _T_265 ? inst[30:25] : _GEN_1840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_1890 = _T_292 ? inst[30:25] : _GEN_1865; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_1915 = _T_321 ? inst[30:25] : _GEN_1890; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] imm_10_5 = io_valid ? _GEN_1915 : 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:62]
  wire [3:0] _GEN_1794 = _T_182 ? inst[11:8] : 4'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:99]
  wire [3:0] _GEN_1819 = _T_209 ? inst[11:8] : _GEN_1794; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] _GEN_1844 = _T_236 ? inst[11:8] : _GEN_1819; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] _GEN_1869 = _T_265 ? inst[11:8] : _GEN_1844; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] _GEN_1894 = _T_292 ? inst[11:8] : _GEN_1869; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] _GEN_1919 = _T_321 ? inst[11:8] : _GEN_1894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] imm_4_1 = io_valid ? _GEN_1919 : 4'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:99]
  wire [12:0] _imm_T_62 = {imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire  imm_signBit_18 = _imm_T_62[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [50:0] _imm_T_64 = imm_signBit_18 ? 51'h7ffffffffffff : 51'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _imm_T_65 = {_imm_T_64,imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  _GEN_1621 = _T_133 & inst[31]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:27]
  wire  imm_20 = io_valid & _GEN_1621; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:27]
  wire [7:0] _GEN_1624 = _T_133 ? inst[19:12] : 8'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:99]
  wire [7:0] imm_19_12 = io_valid ? _GEN_1624 : 8'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:99]
  wire [9:0] _GEN_1622 = _T_133 ? inst[30:21] : 10'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:62]
  wire [9:0] imm_10_1 = io_valid ? _GEN_1622 : 10'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:62]
  wire [20:0] _imm_T_35 = {imm_20,imm_19_12,imm_11,imm_10_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 52:141]
  wire  imm_signBit_11 = _imm_T_35[20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [42:0] _imm_T_37 = imm_signBit_11 ? 43'h7ffffffffff : 43'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _imm_T_38 = {_imm_T_37,imm_20,imm_19_12,imm_11,imm_10_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  _T_59 = 32'h17 == _T_132; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_55 = 32'h37 == _T_132; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _GEN_704 = _T_55 ? inst[31:12] : 20'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 41:27]
  wire [19:0] _GEN_773 = _T_59 ? inst[31:12] : _GEN_704; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [19:0] imm_31_12 = io_valid ? _GEN_773 : 20'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 41:27]
  wire [31:0] _imm_T_31 = {imm_31_12,12'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:141]
  wire  imm_signBit_10 = _imm_T_31[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _imm_T_33 = imm_signBit_10 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _imm_T_34 = {_imm_T_33,imm_31_12,12'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_70 = _T_1 ? _imm_T_321 : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 22:24]
  wire [63:0] _GEN_141 = _T_7 ? _imm_T_321 : _GEN_70; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_212 = _T_13 ? _imm_T_321 : _GEN_141; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_283 = _T_19 ? _imm_T_321 : _GEN_212; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_354 = _T_25 ? _imm_T_321 : _GEN_283; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_425 = _T_31 ? _imm_T_321 : _GEN_354; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_496 = _T_545 ? _imm_T_321 : _GEN_425; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_567 = _T_551 ? _imm_T_321 : _GEN_496; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_638 = _T_557 ? _imm_T_321 : _GEN_567; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_707 = _T_55 ? _imm_T_34 : _GEN_638; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:127]
  wire [63:0] _GEN_776 = _T_59 ? _imm_T_34 : _GEN_707; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:127]
  wire [63:0] _GEN_1627 = _T_133 ? _imm_T_38 : _GEN_776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 52:127]
  wire [63:0] _GEN_1740 = _T_157 ? _imm_T_321 : _GEN_1627; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_1797 = _T_182 ? _imm_T_65 : _GEN_1740; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [63:0] _GEN_1822 = _T_209 ? _imm_T_65 : _GEN_1797; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [63:0] _GEN_1847 = _T_236 ? _imm_T_65 : _GEN_1822; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [63:0] _GEN_1872 = _T_265 ? _imm_T_65 : _GEN_1847; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [63:0] _GEN_1897 = _T_292 ? _imm_T_65 : _GEN_1872; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [63:0] _GEN_1922 = _T_321 ? _imm_T_65 : _GEN_1897; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [63:0] _GEN_2003 = _T_348 ? _imm_T_321 : _GEN_1922; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_2116 = _T_368 ? _imm_T_321 : _GEN_2003; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_2229 = _T_388 ? _imm_T_321 : _GEN_2116; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_2307 = _T_408 ? _imm_T_321 : _GEN_2229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_2420 = _T_427 ? _imm_T_321 : _GEN_2307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_2467 = _T_447 ? _imm_T_132 : _GEN_2420; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:127]
  wire [63:0] _GEN_2487 = _T_470 ? _imm_T_132 : _GEN_2467; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:127]
  wire [63:0] _GEN_2507 = _T_494 ? _imm_T_132 : _GEN_2487; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:127]
  wire [63:0] _GEN_2520 = _T_518 ? _imm_T_321 : _GEN_2507; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_2538 = _T_524 ? _imm_T_321 : _GEN_2520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_2549 = _T_533 ? _imm_T_321 : _GEN_2538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_2588 = _T_539 ? _imm_T_321 : _GEN_2549; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_2659 = _T_545 ? _imm_T_321 : _GEN_2588; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_2730 = _T_551 ? _imm_T_321 : _GEN_2659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_2801 = _T_557 ? _imm_T_321 : _GEN_2730; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_2872 = _T_563 ? _imm_T_321 : _GEN_2801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_2943 = _T_569 ? _imm_T_321 : _GEN_2872; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_3014 = _T_575 ? _imm_T_321 : _GEN_2943; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_3690 = _T_637 ? _imm_T_321 : _GEN_3014; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_3803 = _T_657 ? _imm_T_321 : _GEN_3690; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_3854 = _T_677 ? _imm_T_132 : _GEN_3803; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:127]
  wire [63:0] _GEN_3900 = _T_704 ? _imm_T_141 : _GEN_3854; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 140:20]
  wire [63:0] _GEN_3941 = _T_711 ? _imm_T_150 : _GEN_3900; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 145:11]
  wire [63:0] _GEN_4017 = _T_720 ? _imm_T_166 : _GEN_3941; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 151:28]
  wire [63:0] _GEN_4124 = _T_729 ? _imm_T_166 : _GEN_4017; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 156:11]
  wire [63:0] _GEN_4133 = _T_741 ? _imm_T_198 : _GEN_4124; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 160:21 162:25]
  wire [63:0] _GEN_4202 = _T_770 ? _imm_T_224 : _GEN_4133; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24 188:11]
  wire [63:0] _GEN_4246 = _T_779 ? _imm_T_224 : _GEN_4202; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24 196:11]
  wire [63:0] _GEN_4288 = _T_791 ? _imm_T_309 : _GEN_4246; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22 206:20]
  wire [63:0] _GEN_4611 = _T_862 ? {{58'd0}, _imm_T_306} : _GEN_4288; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24 232:20]
  wire [63:0] _GEN_4715 = _T_875 ? {{58'd0}, _imm_T_306} : _GEN_4611; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24 237:28]
  wire [63:0] _GEN_4819 = _T_889 ? {{58'd0}, _imm_T_306} : _GEN_4715; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24 242:28]
  wire [63:0] _GEN_4923 = _T_897 ? _imm_T_309 : _GEN_4819; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24 247:28]
  wire [63:0] _GEN_5682 = _T_971 ? _imm_T_274 : _GEN_4923; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24 269:20]
  wire [63:0] _GEN_5723 = _T_978 ? _imm_T_283 : _GEN_5682; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24 274:11]
  wire [63:0] _GEN_5799 = _T_987 ? _imm_T_299 : _GEN_5723; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22 280:28]
  wire [63:0] _GEN_5906 = _T_996 ? _imm_T_299 : _GEN_5799; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22 285:11]
  wire [63:0] _GEN_5950 = _T_1011 ? _imm_T_309 : _GEN_5906; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25 292:20]
  wire [63:0] _GEN_7193 = _T_1125 ? _imm_T_321 : _GEN_5950; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [63:0] _GEN_7214 = _T_1132 ? _imm_T_321 : _GEN_7193; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [63:0] _GEN_7228 = _T_1139 ? _imm_T_321 : _GEN_7214; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28]
  wire [63:0] _GEN_7235 = _T_1145 ? _imm_T_321 : _GEN_7228; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28]
  wire [63:0] imm = io_valid ? _GEN_7235 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 22:24]
  wire [63:0] _T_663 = _GEN_31 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:47]
  wire  _T_669 = _T_663[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_667 = _T_663[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_665 = ~_T_663[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire [4:0] _GEN_875 = _T_63 ? inst[24:20] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 20:24]
  wire [4:0] _GEN_946 = _T_70 ? inst[24:20] : _GEN_875; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1017 = _T_77 ? inst[24:20] : _GEN_946; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1088 = _T_84 ? inst[24:20] : _GEN_1017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1159 = _T_91 ? inst[24:20] : _GEN_1088; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1230 = _T_98 ? inst[24:20] : _GEN_1159; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1301 = _T_581 ? inst[24:20] : _GEN_1230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1372 = _T_588 ? inst[24:20] : _GEN_1301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1443 = _T_119 ? inst[24:20] : _GEN_1372; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1514 = _T_595 ? inst[24:20] : _GEN_1443; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1791 = _T_182 ? inst[24:20] : _GEN_1514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1816 = _T_209 ? inst[24:20] : _GEN_1791; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1841 = _T_236 ? inst[24:20] : _GEN_1816; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1866 = _T_265 ? inst[24:20] : _GEN_1841; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1891 = _T_292 ? inst[24:20] : _GEN_1866; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1916 = _T_321 ? inst[24:20] : _GEN_1891; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2462 = _T_447 ? inst[24:20] : _GEN_1916; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2482 = _T_470 ? inst[24:20] : _GEN_2462; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2502 = _T_494 ? inst[24:20] : _GEN_2482; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3081 = _T_581 ? inst[24:20] : _GEN_2502; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3152 = _T_588 ? inst[24:20] : _GEN_3081; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3223 = _T_595 ? inst[24:20] : _GEN_3152; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3294 = _T_602 ? inst[24:20] : _GEN_3223; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3365 = _T_609 ? inst[24:20] : _GEN_3294; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3436 = _T_616 ? inst[24:20] : _GEN_3365; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3507 = _T_623 ? inst[24:20] : _GEN_3436; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3578 = _T_630 ? inst[24:20] : _GEN_3507; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3849 = _T_677 ? inst[24:20] : _GEN_3578; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3939 = _T_711 ? inst[6:2] : _GEN_3849; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4147 = _T_755 ? inst[6:2] : _GEN_3939; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4155 = _T_764 ? inst[6:2] : _GEN_4147; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4991 = _T_911 ? inst[6:2] : _GEN_4155; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5061 = _T_923 ? inst[6:2] : _GEN_4991; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5721 = _T_978 ? inst[6:2] : _GEN_5061; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6287 = _T_1034 ? inst[24:20] : _GEN_5721; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6358 = _T_1041 ? inst[24:20] : _GEN_6287; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6429 = _T_1048 ? inst[24:20] : _GEN_6358; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6500 = _T_1055 ? inst[24:20] : _GEN_6429; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6571 = _T_1062 ? inst[24:20] : _GEN_6500; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6642 = _T_1069 ? inst[24:20] : _GEN_6571; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6713 = _T_1076 ? inst[24:20] : _GEN_6642; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6784 = _T_1083 ? inst[24:20] : _GEN_6713; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6855 = _T_1090 ? inst[24:20] : _GEN_6784; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6926 = _T_1097 ? inst[24:20] : _GEN_6855; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6997 = _T_1104 ? inst[24:20] : _GEN_6926; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7068 = _T_1111 ? inst[24:20] : _GEN_6997; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7139 = _T_1118 ? inst[24:20] : _GEN_7068; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] rs2 = io_valid ? _GEN_7139 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 20:24]
  wire  _GEN_2108 = _T_665 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2152 = _T_368 & _GEN_2108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire  _GEN_2221 = _T_667 ? _GEN_2152 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2265 = _T_388 ? _GEN_2221 : _GEN_2152; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2412 = _T_665 ? _GEN_2265 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2456 = _T_427 ? _GEN_2412 : _GEN_2265; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire  _GEN_3682 = _T_667 ? _GEN_2456 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_3726 = _T_637 ? _GEN_3682 : _GEN_2456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire  _GEN_3795 = _T_669 ? _GEN_3726 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_3839 = _T_657 ? _GEN_3795 : _GEN_3726; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire  exceptionVec_4 = io_valid & _GEN_3839; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_4 = exceptionVec_4 ? 6'h4 : 6'h0; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _GEN_2492 = _T_470 & _GEN_2108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire  _GEN_2498 = _T_667 ? _GEN_2492 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2512 = _T_494 ? _GEN_2498 : _GEN_2492; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire  _GEN_3845 = _T_669 ? _GEN_2512 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_3859 = _T_677 ? _GEN_3845 : _GEN_2512; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire  exceptionVec_6 = io_valid & _GEN_3859; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_5 = exceptionVec_6 ? 6'h6 : _exceptionNO_T_4; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _T_529 = 2'h3 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42]
  wire  _GEN_2527 = 2'h1 == io_now_internal_privilegeMode ? 1'h0 : 2'h0 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_2531 = 2'h3 == io_now_internal_privilegeMode ? 1'h0 : _GEN_2527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_2542 = _T_524 & _GEN_2531; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  exceptionVec_8 = io_valid & _GEN_2542; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_6 = exceptionVec_8 ? 6'h8 : _exceptionNO_T_5; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _GEN_2530 = 2'h3 == io_now_internal_privilegeMode ? 1'h0 : 2'h1 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_2541 = _T_524 & _GEN_2530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  exceptionVec_9 = io_valid & _GEN_2541; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_7 = exceptionVec_9 ? 6'h9 : _exceptionNO_T_6; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _GEN_2539 = _T_524 & _T_529; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  exceptionVec_11 = io_valid & _GEN_2539; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_8 = exceptionVec_11 ? 6'hb : _exceptionNO_T_7; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _GEN_810 = 5'h1 == rs2 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_811 = 5'h2 == rs2 ? io_now_reg_2 : _GEN_810; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_812 = 5'h3 == rs2 ? io_now_reg_3 : _GEN_811; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_813 = 5'h4 == rs2 ? io_now_reg_4 : _GEN_812; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_814 = 5'h5 == rs2 ? io_now_reg_5 : _GEN_813; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_815 = 5'h6 == rs2 ? io_now_reg_6 : _GEN_814; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_816 = 5'h7 == rs2 ? io_now_reg_7 : _GEN_815; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_817 = 5'h8 == rs2 ? io_now_reg_8 : _GEN_816; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_818 = 5'h9 == rs2 ? io_now_reg_9 : _GEN_817; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_819 = 5'ha == rs2 ? io_now_reg_10 : _GEN_818; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_820 = 5'hb == rs2 ? io_now_reg_11 : _GEN_819; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_821 = 5'hc == rs2 ? io_now_reg_12 : _GEN_820; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_822 = 5'hd == rs2 ? io_now_reg_13 : _GEN_821; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_823 = 5'he == rs2 ? io_now_reg_14 : _GEN_822; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_824 = 5'hf == rs2 ? io_now_reg_15 : _GEN_823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_825 = 5'h10 == rs2 ? io_now_reg_16 : _GEN_824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_826 = 5'h11 == rs2 ? io_now_reg_17 : _GEN_825; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_827 = 5'h12 == rs2 ? io_now_reg_18 : _GEN_826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_828 = 5'h13 == rs2 ? io_now_reg_19 : _GEN_827; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_829 = 5'h14 == rs2 ? io_now_reg_20 : _GEN_828; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_830 = 5'h15 == rs2 ? io_now_reg_21 : _GEN_829; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_831 = 5'h16 == rs2 ? io_now_reg_22 : _GEN_830; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_832 = 5'h17 == rs2 ? io_now_reg_23 : _GEN_831; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_833 = 5'h18 == rs2 ? io_now_reg_24 : _GEN_832; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_834 = 5'h19 == rs2 ? io_now_reg_25 : _GEN_833; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_835 = 5'h1a == rs2 ? io_now_reg_26 : _GEN_834; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_836 = 5'h1b == rs2 ? io_now_reg_27 : _GEN_835; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_837 = 5'h1c == rs2 ? io_now_reg_28 : _GEN_836; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_838 = 5'h1d == rs2 ? io_now_reg_29 : _GEN_837; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_839 = 5'h1e == rs2 ? io_now_reg_30 : _GEN_838; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_840 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [1:0] _T_332 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire [63:0] _T_334 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:49]
  wire  _T_340 = _T_334[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_338 = _T_334[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_336 = ~_T_334[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_342 = 2'h1 == _T_332 ? _T_336 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_344 = 2'h2 == _T_332 ? _T_338 : _T_342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_346 = 2'h3 == _T_332 ? _T_340 : _T_344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [63:0] _T_300 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_30; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:25]
  wire [63:0] _T_301 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:48]
  wire  _T_273 = _GEN_31 < _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:25]
  wire  _T_246 = $signed(_T_300) < $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:32]
  wire [63:0] _T_168 = {_T_663[63:1],1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:43]
  wire  _T_174 = _T_168[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_172 = _T_168[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_170 = ~_T_168[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_176 = 2'h1 == _T_332 ? _T_170 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_178 = 2'h2 == _T_332 ? _T_172 : _T_176; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_180 = 2'h3 == _T_332 ? _T_174 : _T_178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _GEN_1618 = _T_346 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30 144:33]
  wire  _GEN_1663 = _T_133 & _GEN_1618; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_1732 = _T_180 ? _GEN_1663 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1776 = _T_157 ? _GEN_1732 : _GEN_1663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire  _GEN_1781 = _T_346 ? _GEN_1776 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1786 = _GEN_31 == _GEN_840 ? _GEN_1781 : _GEN_1776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire  _GEN_1801 = _T_182 ? _GEN_1786 : _GEN_1776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire  _GEN_1806 = _T_346 ? _GEN_1801 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1811 = _GEN_31 != _GEN_840 ? _GEN_1806 : _GEN_1801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire  _GEN_1826 = _T_209 ? _GEN_1811 : _GEN_1801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire  _GEN_1831 = _T_346 ? _GEN_1826 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1836 = $signed(_T_300) < $signed(_T_301) ? _GEN_1831 : _GEN_1826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire  _GEN_1851 = _T_236 ? _GEN_1836 : _GEN_1826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire  _GEN_1856 = _T_346 ? _GEN_1851 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1861 = _GEN_31 < _GEN_840 ? _GEN_1856 : _GEN_1851; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire  _GEN_1876 = _T_265 ? _GEN_1861 : _GEN_1851; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire  _GEN_1881 = _T_346 ? _GEN_1876 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1886 = $signed(_T_300) >= $signed(_T_301) ? _GEN_1881 : _GEN_1876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire  _GEN_1901 = _T_292 ? _GEN_1886 : _GEN_1876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire  _GEN_1906 = _T_346 ? _GEN_1901 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1911 = _GEN_31 >= _GEN_840 ? _GEN_1906 : _GEN_1901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire  _GEN_1926 = _T_321 ? _GEN_1911 : _GEN_1901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire  exceptionVec_0 = io_valid & _GEN_1926; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_9 = exceptionVec_0 ? 6'h0 : _exceptionNO_T_8; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _T_1025 = inst & 32'hfc63; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1026 = 32'h9c01 == _T_1025; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1018 = 32'h9c21 == _T_1025; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_953 = 32'h8c01 == _T_1025; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_945 = 32'h8c21 == _T_1025; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_937 = 32'h8c41 == _T_1025; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_929 = 32'h8c61 == _T_1025; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_845 = inst[12:5] != 8'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 23:96]
  wire  _T_846 = 32'h0 == _T_1007 & _T_845; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _GEN_64 = _T_1 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 125:24 128:24]
  wire  _GEN_135 = _T_7 ? 1'h0 : _GEN_64; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_206 = _T_13 ? 1'h0 : _GEN_135; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_277 = _T_19 ? 1'h0 : _GEN_206; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_348 = _T_25 ? 1'h0 : _GEN_277; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_419 = _T_31 ? 1'h0 : _GEN_348; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_490 = _T_545 ? 1'h0 : _GEN_419; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_561 = _T_551 ? 1'h0 : _GEN_490; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_632 = _T_557 ? 1'h0 : _GEN_561; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_703 = _T_55 ? 1'h0 : _GEN_632; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_772 = _T_59 ? 1'h0 : _GEN_703; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_873 = _T_63 ? 1'h0 : _GEN_772; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_944 = _T_70 ? 1'h0 : _GEN_873; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1015 = _T_77 ? 1'h0 : _GEN_944; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1086 = _T_84 ? 1'h0 : _GEN_1015; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1157 = _T_91 ? 1'h0 : _GEN_1086; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1228 = _T_98 ? 1'h0 : _GEN_1157; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1299 = _T_581 ? 1'h0 : _GEN_1228; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1370 = _T_588 ? 1'h0 : _GEN_1299; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1441 = _T_119 ? 1'h0 : _GEN_1370; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1512 = _T_595 ? 1'h0 : _GEN_1441; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1620 = _T_133 ? 1'h0 : _GEN_1512; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1734 = _T_157 ? 1'h0 : _GEN_1620; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1788 = _T_182 ? 1'h0 : _GEN_1734; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1813 = _T_209 ? 1'h0 : _GEN_1788; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1838 = _T_236 ? 1'h0 : _GEN_1813; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1863 = _T_265 ? 1'h0 : _GEN_1838; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1888 = _T_292 ? 1'h0 : _GEN_1863; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1913 = _T_321 ? 1'h0 : _GEN_1888; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1997 = _T_348 ? 1'h0 : _GEN_1913; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2110 = _T_368 ? 1'h0 : _GEN_1997; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2223 = _T_388 ? 1'h0 : _GEN_2110; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2301 = _T_408 ? 1'h0 : _GEN_2223; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2414 = _T_427 ? 1'h0 : _GEN_2301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2460 = _T_447 ? 1'h0 : _GEN_2414; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2480 = _T_470 ? 1'h0 : _GEN_2460; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2500 = _T_494 ? 1'h0 : _GEN_2480; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2514 = _T_518 ? 1'h0 : _GEN_2500; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2532 = _T_524 ? 1'h0 : _GEN_2514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2543 = _T_533 ? 1'h0 : _GEN_2532; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2582 = _T_539 ? 1'h0 : _GEN_2543; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2653 = _T_545 ? 1'h0 : _GEN_2582; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2724 = _T_551 ? 1'h0 : _GEN_2653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2795 = _T_557 ? 1'h0 : _GEN_2724; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2866 = _T_563 ? 1'h0 : _GEN_2795; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2937 = _T_569 ? 1'h0 : _GEN_2866; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3008 = _T_575 ? 1'h0 : _GEN_2937; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3079 = _T_581 ? 1'h0 : _GEN_3008; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3150 = _T_588 ? 1'h0 : _GEN_3079; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3221 = _T_595 ? 1'h0 : _GEN_3150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3292 = _T_602 ? 1'h0 : _GEN_3221; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3363 = _T_609 ? 1'h0 : _GEN_3292; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3434 = _T_616 ? 1'h0 : _GEN_3363; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3505 = _T_623 ? 1'h0 : _GEN_3434; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3576 = _T_630 ? 1'h0 : _GEN_3505; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3684 = _T_637 ? 1'h0 : _GEN_3576; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3797 = _T_657 ? 1'h0 : _GEN_3684; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3847 = _T_677 ? 1'h0 : _GEN_3797; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3893 = _T_704 ? 1'h0 : _GEN_3847; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3936 = _T_711 ? 1'h0 : _GEN_3893; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4010 = _T_720 ? 1'h0 : _GEN_3936; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4117 = _T_729 ? 1'h0 : _GEN_4010; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4129 = _T_741 ? 1'h0 : _GEN_4117; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 160:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4144 = _T_755 ? 1'h0 : _GEN_4129; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4152 = _T_764 ? 1'h0 : _GEN_4144; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4195 = _T_770 ? 1'h0 : _GEN_4152; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4239 = _T_779 ? 1'h0 : _GEN_4195; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4281 = _T_791 ? 1'h0 : _GEN_4239; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4353 = _T_809 ? 1'h0 : _GEN_4281; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4456 = _T_824 ? 1'h0 : _GEN_4353; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4495 = _T_836 ? 1'h0 : _GEN_4456; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 220:28 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4535 = _T_846 ? 1'h0 : _GEN_4495; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4604 = _T_862 ? 1'h0 : _GEN_4535; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4708 = _T_875 ? 1'h0 : _GEN_4604; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4812 = _T_889 ? 1'h0 : _GEN_4708; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4916 = _T_897 ? 1'h0 : _GEN_4812; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4988 = _T_911 ? 1'h0 : _GEN_4916; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5058 = _T_923 ? 1'h0 : _GEN_4988; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5192 = _T_929 ? 1'h0 : _GEN_5058; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5327 = _T_937 ? 1'h0 : _GEN_5192; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5462 = _T_945 ? 1'h0 : _GEN_5327; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5597 = _T_953 ? 1'h0 : _GEN_5462; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5636 = _T_961 ? 1'h0 : _GEN_5597; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 259:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5675 = _T_971 ? 1'h0 : _GEN_5636; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5718 = _T_978 ? 1'h0 : _GEN_5675; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5792 = _T_987 ? 1'h0 : _GEN_5718; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5899 = _T_996 ? 1'h0 : _GEN_5792; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5943 = _T_1011 ? 1'h0 : _GEN_5899; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6079 = _T_1018 ? 1'h0 : _GEN_5943; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6214 = _T_1026 ? 1'h0 : _GEN_6079; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6285 = _T_1034 ? 1'h0 : _GEN_6214; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6356 = _T_1041 ? 1'h0 : _GEN_6285; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6427 = _T_1048 ? 1'h0 : _GEN_6356; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6498 = _T_1055 ? 1'h0 : _GEN_6427; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6569 = _T_1062 ? 1'h0 : _GEN_6498; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6640 = _T_1069 ? 1'h0 : _GEN_6569; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6711 = _T_1076 ? 1'h0 : _GEN_6640; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6782 = _T_1083 ? 1'h0 : _GEN_6711; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6853 = _T_1090 ? 1'h0 : _GEN_6782; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6924 = _T_1097 ? 1'h0 : _GEN_6853; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6995 = _T_1104 ? 1'h0 : _GEN_6924; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_7066 = _T_1111 ? 1'h0 : _GEN_6995; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_7137 = _T_1118 ? 1'h0 : _GEN_7066; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_7187 = _T_1125 ? 1'h0 : _GEN_7137; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_7208 = _T_1132 ? 1'h0 : _GEN_7187; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_7222 = _T_1139 ? 1'h0 : _GEN_7208; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_7229 = _T_1145 ? 1'h0 : _GEN_7222; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  illegalInstruction = io_valid & _GEN_7229; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 119:36]
  wire  illegalSret = io_now_internal_privilegeMode < 2'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 118:55]
  wire  mstatusOld_tsr = io_now_csr_mstatus[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  illegalSModeSret = io_now_internal_privilegeMode == 2'h1 & mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 119:65]
  wire  _T_1130 = illegalSret | illegalSModeSret; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:22]
  wire  _GEN_7194 = _T_1125 & _T_1130; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_7206 = io_now_internal_privilegeMode == 2'h3 ? _GEN_7194 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 88:48 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_7220 = _T_1132 ? _GEN_7206 : _GEN_7194; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire  _GEN_7237 = illegalInstruction | _GEN_7220; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 133:30 144:33]
  wire  exceptionVec_2 = io_valid & _GEN_7237; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_10 = exceptionVec_2 ? 6'h2 : _exceptionNO_T_9; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  exceptionVec_3 = io_valid & _T_518; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] exceptionNO = exceptionVec_3 ? 6'h3 : _exceptionNO_T_10; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [4:0] _GEN_68 = _T_1 ? inst[11:7] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 17:24]
  wire [4:0] _GEN_139 = _T_7 ? inst[11:7] : _GEN_68; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_210 = _T_13 ? inst[11:7] : _GEN_139; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_281 = _T_19 ? inst[11:7] : _GEN_210; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_352 = _T_25 ? inst[11:7] : _GEN_281; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_423 = _T_31 ? inst[11:7] : _GEN_352; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_494 = _T_545 ? inst[11:7] : _GEN_423; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_565 = _T_551 ? inst[11:7] : _GEN_494; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_636 = _T_557 ? inst[11:7] : _GEN_565; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_705 = _T_55 ? inst[11:7] : _GEN_636; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_774 = _T_59 ? inst[11:7] : _GEN_705; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_878 = _T_63 ? inst[11:7] : _GEN_774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_949 = _T_70 ? inst[11:7] : _GEN_878; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1020 = _T_77 ? inst[11:7] : _GEN_949; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1091 = _T_84 ? inst[11:7] : _GEN_1020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1162 = _T_91 ? inst[11:7] : _GEN_1091; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1233 = _T_98 ? inst[11:7] : _GEN_1162; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1304 = _T_581 ? inst[11:7] : _GEN_1233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1375 = _T_588 ? inst[11:7] : _GEN_1304; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1446 = _T_119 ? inst[11:7] : _GEN_1375; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1517 = _T_595 ? inst[11:7] : _GEN_1446; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1625 = _T_133 ? inst[11:7] : _GEN_1517; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1738 = _T_157 ? inst[11:7] : _GEN_1625; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2001 = _T_348 ? inst[11:7] : _GEN_1738; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2114 = _T_368 ? inst[11:7] : _GEN_2001; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2227 = _T_388 ? inst[11:7] : _GEN_2114; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2305 = _T_408 ? inst[11:7] : _GEN_2227; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2418 = _T_427 ? inst[11:7] : _GEN_2305; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2518 = _T_518 ? inst[11:7] : _GEN_2418; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2536 = _T_524 ? inst[11:7] : _GEN_2518; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2547 = _T_533 ? inst[11:7] : _GEN_2536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2586 = _T_539 ? inst[11:7] : _GEN_2547; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2657 = _T_545 ? inst[11:7] : _GEN_2586; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2728 = _T_551 ? inst[11:7] : _GEN_2657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2799 = _T_557 ? inst[11:7] : _GEN_2728; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2870 = _T_563 ? inst[11:7] : _GEN_2799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2941 = _T_569 ? inst[11:7] : _GEN_2870; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3012 = _T_575 ? inst[11:7] : _GEN_2941; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3084 = _T_581 ? inst[11:7] : _GEN_3012; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3155 = _T_588 ? inst[11:7] : _GEN_3084; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3226 = _T_595 ? inst[11:7] : _GEN_3155; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3297 = _T_602 ? inst[11:7] : _GEN_3226; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3368 = _T_609 ? inst[11:7] : _GEN_3297; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3439 = _T_616 ? inst[11:7] : _GEN_3368; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3510 = _T_623 ? inst[11:7] : _GEN_3439; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3581 = _T_630 ? inst[11:7] : _GEN_3510; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3688 = _T_637 ? inst[11:7] : _GEN_3581; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3801 = _T_657 ? inst[11:7] : _GEN_3688; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3899 = _T_704 ? rs1 : _GEN_3801; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 138:24]
  wire [4:0] _GEN_4149 = _T_755 ? rs1 : _GEN_3899; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 112:110 173:22]
  wire [4:0] _GEN_4157 = _T_764 ? rs1 : _GEN_4149; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 112:110 179:24]
  wire [4:0] _GEN_4287 = _T_791 ? rs1 : _GEN_4157; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 204:22]
  wire [4:0] _GEN_4359 = _T_809 ? rs1 : _GEN_4287; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 209:23]
  wire [4:0] _GEN_4462 = _T_824 ? rs1 : _GEN_4359; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 215:24]
  wire [4:0] _GEN_4501 = _T_836 ? rs1 : _GEN_4462; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 220:28]
  wire [4:0] _GEN_4610 = _T_862 ? rs1 : _GEN_4501; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 230:24]
  wire [4:0] _GEN_4993 = _T_911 ? rs1 : _GEN_4610; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 112:110 251:23]
  wire [4:0] _GEN_5063 = _T_923 ? rs1 : _GEN_4993; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 112:110 252:23]
  wire [4:0] _GEN_5642 = _T_961 ? rs1 : _GEN_5063; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 259:23]
  wire [4:0] _GEN_5681 = _T_971 ? rs1 : _GEN_5642; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 267:24]
  wire [4:0] _GEN_5949 = _T_1011 ? rs1 : _GEN_5681; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 290:25]
  wire [4:0] _GEN_6290 = _T_1034 ? inst[11:7] : _GEN_5949; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6361 = _T_1041 ? inst[11:7] : _GEN_6290; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6432 = _T_1048 ? inst[11:7] : _GEN_6361; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6503 = _T_1055 ? inst[11:7] : _GEN_6432; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6574 = _T_1062 ? inst[11:7] : _GEN_6503; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6645 = _T_1069 ? inst[11:7] : _GEN_6574; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6716 = _T_1076 ? inst[11:7] : _GEN_6645; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6787 = _T_1083 ? inst[11:7] : _GEN_6716; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6858 = _T_1090 ? inst[11:7] : _GEN_6787; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6929 = _T_1097 ? inst[11:7] : _GEN_6858; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7000 = _T_1104 ? inst[11:7] : _GEN_6929; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7071 = _T_1111 ? inst[11:7] : _GEN_7000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7142 = _T_1118 ? inst[11:7] : _GEN_7071; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7191 = _T_1125 ? inst[11:7] : _GEN_7142; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7212 = _T_1132 ? inst[11:7] : _GEN_7191; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7226 = _T_1139 ? inst[11:7] : _GEN_7212; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7233 = _T_1145 ? inst[11:7] : _GEN_7226; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] rd = io_valid ? _GEN_7233 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 17:24]
  wire [63:0] _GEN_33 = 5'h1 == rd ? _T_663 : io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_34 = 5'h2 == rd ? _T_663 : io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_35 = 5'h3 == rd ? _T_663 : io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_36 = 5'h4 == rd ? _T_663 : io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_37 = 5'h5 == rd ? _T_663 : io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_38 = 5'h6 == rd ? _T_663 : io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_39 = 5'h7 == rd ? _T_663 : io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_40 = 5'h8 == rd ? _T_663 : io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_41 = 5'h9 == rd ? _T_663 : io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_42 = 5'ha == rd ? _T_663 : io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_43 = 5'hb == rd ? _T_663 : io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_44 = 5'hc == rd ? _T_663 : io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_45 = 5'hd == rd ? _T_663 : io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_46 = 5'he == rd ? _T_663 : io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_47 = 5'hf == rd ? _T_663 : io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_48 = 5'h10 == rd ? _T_663 : io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_49 = 5'h11 == rd ? _T_663 : io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_50 = 5'h12 == rd ? _T_663 : io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_51 = 5'h13 == rd ? _T_663 : io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_52 = 5'h14 == rd ? _T_663 : io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_53 = 5'h15 == rd ? _T_663 : io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_54 = 5'h16 == rd ? _T_663 : io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_55 = 5'h17 == rd ? _T_663 : io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_56 = 5'h18 == rd ? _T_663 : io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_57 = 5'h19 == rd ? _T_663 : io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_58 = 5'h1a == rd ? _T_663 : io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_59 = 5'h1b == rd ? _T_663 : io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_60 = 5'h1c == rd ? _T_663 : io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_61 = 5'h1d == rd ? _T_663 : io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_62 = 5'h1e == rd ? _T_663 : io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_63 = 5'h1f == rd ? _T_663 : io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_72 = _T_1 ? _GEN_33 : io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_73 = _T_1 ? _GEN_34 : io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_74 = _T_1 ? _GEN_35 : io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_75 = _T_1 ? _GEN_36 : io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_76 = _T_1 ? _GEN_37 : io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_77 = _T_1 ? _GEN_38 : io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_78 = _T_1 ? _GEN_39 : io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_79 = _T_1 ? _GEN_40 : io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_80 = _T_1 ? _GEN_41 : io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_81 = _T_1 ? _GEN_42 : io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_82 = _T_1 ? _GEN_43 : io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_83 = _T_1 ? _GEN_44 : io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_84 = _T_1 ? _GEN_45 : io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_85 = _T_1 ? _GEN_46 : io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_86 = _T_1 ? _GEN_47 : io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_87 = _T_1 ? _GEN_48 : io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_88 = _T_1 ? _GEN_49 : io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_89 = _T_1 ? _GEN_50 : io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_90 = _T_1 ? _GEN_51 : io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_91 = _T_1 ? _GEN_52 : io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_92 = _T_1 ? _GEN_53 : io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_93 = _T_1 ? _GEN_54 : io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_94 = _T_1 ? _GEN_55 : io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_95 = _T_1 ? _GEN_56 : io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_96 = _T_1 ? _GEN_57 : io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_97 = _T_1 ? _GEN_58 : io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_98 = _T_1 ? _GEN_59 : io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_99 = _T_1 ? _GEN_60 : io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_100 = _T_1 ? _GEN_61 : io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_101 = _T_1 ? _GEN_62 : io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_102 = _T_1 ? _GEN_63 : io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _next_reg_T_3 = io_valid ? _GEN_7235 : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:80]
  wire [63:0] _next_reg_rd_0 = {{63'd0}, $signed(_T_300) < $signed(_next_reg_T_3)}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_104 = 5'h1 == rd ? _next_reg_rd_0 : _GEN_72; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_105 = 5'h2 == rd ? _next_reg_rd_0 : _GEN_73; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_106 = 5'h3 == rd ? _next_reg_rd_0 : _GEN_74; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_107 = 5'h4 == rd ? _next_reg_rd_0 : _GEN_75; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_108 = 5'h5 == rd ? _next_reg_rd_0 : _GEN_76; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_109 = 5'h6 == rd ? _next_reg_rd_0 : _GEN_77; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_110 = 5'h7 == rd ? _next_reg_rd_0 : _GEN_78; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_111 = 5'h8 == rd ? _next_reg_rd_0 : _GEN_79; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_112 = 5'h9 == rd ? _next_reg_rd_0 : _GEN_80; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_113 = 5'ha == rd ? _next_reg_rd_0 : _GEN_81; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_114 = 5'hb == rd ? _next_reg_rd_0 : _GEN_82; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_115 = 5'hc == rd ? _next_reg_rd_0 : _GEN_83; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_116 = 5'hd == rd ? _next_reg_rd_0 : _GEN_84; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_117 = 5'he == rd ? _next_reg_rd_0 : _GEN_85; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_118 = 5'hf == rd ? _next_reg_rd_0 : _GEN_86; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_119 = 5'h10 == rd ? _next_reg_rd_0 : _GEN_87; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_120 = 5'h11 == rd ? _next_reg_rd_0 : _GEN_88; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_121 = 5'h12 == rd ? _next_reg_rd_0 : _GEN_89; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_122 = 5'h13 == rd ? _next_reg_rd_0 : _GEN_90; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_123 = 5'h14 == rd ? _next_reg_rd_0 : _GEN_91; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_124 = 5'h15 == rd ? _next_reg_rd_0 : _GEN_92; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_125 = 5'h16 == rd ? _next_reg_rd_0 : _GEN_93; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_126 = 5'h17 == rd ? _next_reg_rd_0 : _GEN_94; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_127 = 5'h18 == rd ? _next_reg_rd_0 : _GEN_95; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_128 = 5'h19 == rd ? _next_reg_rd_0 : _GEN_96; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_129 = 5'h1a == rd ? _next_reg_rd_0 : _GEN_97; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_130 = 5'h1b == rd ? _next_reg_rd_0 : _GEN_98; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_131 = 5'h1c == rd ? _next_reg_rd_0 : _GEN_99; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_132 = 5'h1d == rd ? _next_reg_rd_0 : _GEN_100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_133 = 5'h1e == rd ? _next_reg_rd_0 : _GEN_101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_134 = 5'h1f == rd ? _next_reg_rd_0 : _GEN_102; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_143 = _T_7 ? _GEN_104 : _GEN_72; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_144 = _T_7 ? _GEN_105 : _GEN_73; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_145 = _T_7 ? _GEN_106 : _GEN_74; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_146 = _T_7 ? _GEN_107 : _GEN_75; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_147 = _T_7 ? _GEN_108 : _GEN_76; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_148 = _T_7 ? _GEN_109 : _GEN_77; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_149 = _T_7 ? _GEN_110 : _GEN_78; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_150 = _T_7 ? _GEN_111 : _GEN_79; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_151 = _T_7 ? _GEN_112 : _GEN_80; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_152 = _T_7 ? _GEN_113 : _GEN_81; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_153 = _T_7 ? _GEN_114 : _GEN_82; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_154 = _T_7 ? _GEN_115 : _GEN_83; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_155 = _T_7 ? _GEN_116 : _GEN_84; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_156 = _T_7 ? _GEN_117 : _GEN_85; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_157 = _T_7 ? _GEN_118 : _GEN_86; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_158 = _T_7 ? _GEN_119 : _GEN_87; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_159 = _T_7 ? _GEN_120 : _GEN_88; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_160 = _T_7 ? _GEN_121 : _GEN_89; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_161 = _T_7 ? _GEN_122 : _GEN_90; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_162 = _T_7 ? _GEN_123 : _GEN_91; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_163 = _T_7 ? _GEN_124 : _GEN_92; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_164 = _T_7 ? _GEN_125 : _GEN_93; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_165 = _T_7 ? _GEN_126 : _GEN_94; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_166 = _T_7 ? _GEN_127 : _GEN_95; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_167 = _T_7 ? _GEN_128 : _GEN_96; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_168 = _T_7 ? _GEN_129 : _GEN_97; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_169 = _T_7 ? _GEN_130 : _GEN_98; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_170 = _T_7 ? _GEN_131 : _GEN_99; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_171 = _T_7 ? _GEN_132 : _GEN_100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_172 = _T_7 ? _GEN_133 : _GEN_101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_173 = _T_7 ? _GEN_134 : _GEN_102; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _next_reg_rd_1 = {{63'd0}, _GEN_31 < imm}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_175 = 5'h1 == rd ? _next_reg_rd_1 : _GEN_143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_176 = 5'h2 == rd ? _next_reg_rd_1 : _GEN_144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_177 = 5'h3 == rd ? _next_reg_rd_1 : _GEN_145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_178 = 5'h4 == rd ? _next_reg_rd_1 : _GEN_146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_179 = 5'h5 == rd ? _next_reg_rd_1 : _GEN_147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_180 = 5'h6 == rd ? _next_reg_rd_1 : _GEN_148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_181 = 5'h7 == rd ? _next_reg_rd_1 : _GEN_149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_182 = 5'h8 == rd ? _next_reg_rd_1 : _GEN_150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_183 = 5'h9 == rd ? _next_reg_rd_1 : _GEN_151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_184 = 5'ha == rd ? _next_reg_rd_1 : _GEN_152; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_185 = 5'hb == rd ? _next_reg_rd_1 : _GEN_153; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_186 = 5'hc == rd ? _next_reg_rd_1 : _GEN_154; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_187 = 5'hd == rd ? _next_reg_rd_1 : _GEN_155; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_188 = 5'he == rd ? _next_reg_rd_1 : _GEN_156; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_189 = 5'hf == rd ? _next_reg_rd_1 : _GEN_157; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_190 = 5'h10 == rd ? _next_reg_rd_1 : _GEN_158; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_191 = 5'h11 == rd ? _next_reg_rd_1 : _GEN_159; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_192 = 5'h12 == rd ? _next_reg_rd_1 : _GEN_160; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_193 = 5'h13 == rd ? _next_reg_rd_1 : _GEN_161; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_194 = 5'h14 == rd ? _next_reg_rd_1 : _GEN_162; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_195 = 5'h15 == rd ? _next_reg_rd_1 : _GEN_163; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_196 = 5'h16 == rd ? _next_reg_rd_1 : _GEN_164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_197 = 5'h17 == rd ? _next_reg_rd_1 : _GEN_165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_198 = 5'h18 == rd ? _next_reg_rd_1 : _GEN_166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_199 = 5'h19 == rd ? _next_reg_rd_1 : _GEN_167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_200 = 5'h1a == rd ? _next_reg_rd_1 : _GEN_168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_201 = 5'h1b == rd ? _next_reg_rd_1 : _GEN_169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_202 = 5'h1c == rd ? _next_reg_rd_1 : _GEN_170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_203 = 5'h1d == rd ? _next_reg_rd_1 : _GEN_171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_204 = 5'h1e == rd ? _next_reg_rd_1 : _GEN_172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_205 = 5'h1f == rd ? _next_reg_rd_1 : _GEN_173; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_214 = _T_13 ? _GEN_175 : _GEN_143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_215 = _T_13 ? _GEN_176 : _GEN_144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_216 = _T_13 ? _GEN_177 : _GEN_145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_217 = _T_13 ? _GEN_178 : _GEN_146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_218 = _T_13 ? _GEN_179 : _GEN_147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_219 = _T_13 ? _GEN_180 : _GEN_148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_220 = _T_13 ? _GEN_181 : _GEN_149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_221 = _T_13 ? _GEN_182 : _GEN_150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_222 = _T_13 ? _GEN_183 : _GEN_151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_223 = _T_13 ? _GEN_184 : _GEN_152; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_224 = _T_13 ? _GEN_185 : _GEN_153; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_225 = _T_13 ? _GEN_186 : _GEN_154; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_226 = _T_13 ? _GEN_187 : _GEN_155; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_227 = _T_13 ? _GEN_188 : _GEN_156; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_228 = _T_13 ? _GEN_189 : _GEN_157; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_229 = _T_13 ? _GEN_190 : _GEN_158; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_230 = _T_13 ? _GEN_191 : _GEN_159; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_231 = _T_13 ? _GEN_192 : _GEN_160; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_232 = _T_13 ? _GEN_193 : _GEN_161; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_233 = _T_13 ? _GEN_194 : _GEN_162; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_234 = _T_13 ? _GEN_195 : _GEN_163; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_235 = _T_13 ? _GEN_196 : _GEN_164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_236 = _T_13 ? _GEN_197 : _GEN_165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_237 = _T_13 ? _GEN_198 : _GEN_166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_238 = _T_13 ? _GEN_199 : _GEN_167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_239 = _T_13 ? _GEN_200 : _GEN_168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_240 = _T_13 ? _GEN_201 : _GEN_169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_241 = _T_13 ? _GEN_202 : _GEN_170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_242 = _T_13 ? _GEN_203 : _GEN_171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_243 = _T_13 ? _GEN_204 : _GEN_172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_244 = _T_13 ? _GEN_205 : _GEN_173; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _next_reg_T_8 = _GEN_31 & imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:62]
  wire [63:0] _GEN_246 = 5'h1 == rd ? _next_reg_T_8 : _GEN_214; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_247 = 5'h2 == rd ? _next_reg_T_8 : _GEN_215; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_248 = 5'h3 == rd ? _next_reg_T_8 : _GEN_216; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_249 = 5'h4 == rd ? _next_reg_T_8 : _GEN_217; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_250 = 5'h5 == rd ? _next_reg_T_8 : _GEN_218; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_251 = 5'h6 == rd ? _next_reg_T_8 : _GEN_219; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_252 = 5'h7 == rd ? _next_reg_T_8 : _GEN_220; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_253 = 5'h8 == rd ? _next_reg_T_8 : _GEN_221; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_254 = 5'h9 == rd ? _next_reg_T_8 : _GEN_222; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_255 = 5'ha == rd ? _next_reg_T_8 : _GEN_223; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_256 = 5'hb == rd ? _next_reg_T_8 : _GEN_224; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_257 = 5'hc == rd ? _next_reg_T_8 : _GEN_225; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_258 = 5'hd == rd ? _next_reg_T_8 : _GEN_226; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_259 = 5'he == rd ? _next_reg_T_8 : _GEN_227; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_260 = 5'hf == rd ? _next_reg_T_8 : _GEN_228; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_261 = 5'h10 == rd ? _next_reg_T_8 : _GEN_229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_262 = 5'h11 == rd ? _next_reg_T_8 : _GEN_230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_263 = 5'h12 == rd ? _next_reg_T_8 : _GEN_231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_264 = 5'h13 == rd ? _next_reg_T_8 : _GEN_232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_265 = 5'h14 == rd ? _next_reg_T_8 : _GEN_233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_266 = 5'h15 == rd ? _next_reg_T_8 : _GEN_234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_267 = 5'h16 == rd ? _next_reg_T_8 : _GEN_235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_268 = 5'h17 == rd ? _next_reg_T_8 : _GEN_236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_269 = 5'h18 == rd ? _next_reg_T_8 : _GEN_237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_270 = 5'h19 == rd ? _next_reg_T_8 : _GEN_238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_271 = 5'h1a == rd ? _next_reg_T_8 : _GEN_239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_272 = 5'h1b == rd ? _next_reg_T_8 : _GEN_240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_273 = 5'h1c == rd ? _next_reg_T_8 : _GEN_241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_274 = 5'h1d == rd ? _next_reg_T_8 : _GEN_242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_275 = 5'h1e == rd ? _next_reg_T_8 : _GEN_243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_276 = 5'h1f == rd ? _next_reg_T_8 : _GEN_244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_285 = _T_19 ? _GEN_246 : _GEN_214; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_286 = _T_19 ? _GEN_247 : _GEN_215; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_287 = _T_19 ? _GEN_248 : _GEN_216; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_288 = _T_19 ? _GEN_249 : _GEN_217; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_289 = _T_19 ? _GEN_250 : _GEN_218; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_290 = _T_19 ? _GEN_251 : _GEN_219; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_291 = _T_19 ? _GEN_252 : _GEN_220; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_292 = _T_19 ? _GEN_253 : _GEN_221; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_293 = _T_19 ? _GEN_254 : _GEN_222; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_294 = _T_19 ? _GEN_255 : _GEN_223; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_295 = _T_19 ? _GEN_256 : _GEN_224; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_296 = _T_19 ? _GEN_257 : _GEN_225; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_297 = _T_19 ? _GEN_258 : _GEN_226; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_298 = _T_19 ? _GEN_259 : _GEN_227; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_299 = _T_19 ? _GEN_260 : _GEN_228; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_300 = _T_19 ? _GEN_261 : _GEN_229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_301 = _T_19 ? _GEN_262 : _GEN_230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_302 = _T_19 ? _GEN_263 : _GEN_231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_303 = _T_19 ? _GEN_264 : _GEN_232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_304 = _T_19 ? _GEN_265 : _GEN_233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_305 = _T_19 ? _GEN_266 : _GEN_234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_306 = _T_19 ? _GEN_267 : _GEN_235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_307 = _T_19 ? _GEN_268 : _GEN_236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_308 = _T_19 ? _GEN_269 : _GEN_237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_309 = _T_19 ? _GEN_270 : _GEN_238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_310 = _T_19 ? _GEN_271 : _GEN_239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_311 = _T_19 ? _GEN_272 : _GEN_240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_312 = _T_19 ? _GEN_273 : _GEN_241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_313 = _T_19 ? _GEN_274 : _GEN_242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_314 = _T_19 ? _GEN_275 : _GEN_243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_315 = _T_19 ? _GEN_276 : _GEN_244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _next_reg_T_9 = _GEN_31 | imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:62]
  wire [63:0] _GEN_317 = 5'h1 == rd ? _next_reg_T_9 : _GEN_285; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_318 = 5'h2 == rd ? _next_reg_T_9 : _GEN_286; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_319 = 5'h3 == rd ? _next_reg_T_9 : _GEN_287; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_320 = 5'h4 == rd ? _next_reg_T_9 : _GEN_288; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_321 = 5'h5 == rd ? _next_reg_T_9 : _GEN_289; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_322 = 5'h6 == rd ? _next_reg_T_9 : _GEN_290; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_323 = 5'h7 == rd ? _next_reg_T_9 : _GEN_291; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_324 = 5'h8 == rd ? _next_reg_T_9 : _GEN_292; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_325 = 5'h9 == rd ? _next_reg_T_9 : _GEN_293; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_326 = 5'ha == rd ? _next_reg_T_9 : _GEN_294; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_327 = 5'hb == rd ? _next_reg_T_9 : _GEN_295; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_328 = 5'hc == rd ? _next_reg_T_9 : _GEN_296; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_329 = 5'hd == rd ? _next_reg_T_9 : _GEN_297; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_330 = 5'he == rd ? _next_reg_T_9 : _GEN_298; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_331 = 5'hf == rd ? _next_reg_T_9 : _GEN_299; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_332 = 5'h10 == rd ? _next_reg_T_9 : _GEN_300; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_333 = 5'h11 == rd ? _next_reg_T_9 : _GEN_301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_334 = 5'h12 == rd ? _next_reg_T_9 : _GEN_302; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_335 = 5'h13 == rd ? _next_reg_T_9 : _GEN_303; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_336 = 5'h14 == rd ? _next_reg_T_9 : _GEN_304; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_337 = 5'h15 == rd ? _next_reg_T_9 : _GEN_305; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_338 = 5'h16 == rd ? _next_reg_T_9 : _GEN_306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_339 = 5'h17 == rd ? _next_reg_T_9 : _GEN_307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_340 = 5'h18 == rd ? _next_reg_T_9 : _GEN_308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_341 = 5'h19 == rd ? _next_reg_T_9 : _GEN_309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_342 = 5'h1a == rd ? _next_reg_T_9 : _GEN_310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_343 = 5'h1b == rd ? _next_reg_T_9 : _GEN_311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_344 = 5'h1c == rd ? _next_reg_T_9 : _GEN_312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_345 = 5'h1d == rd ? _next_reg_T_9 : _GEN_313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_346 = 5'h1e == rd ? _next_reg_T_9 : _GEN_314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_347 = 5'h1f == rd ? _next_reg_T_9 : _GEN_315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_356 = _T_25 ? _GEN_317 : _GEN_285; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_357 = _T_25 ? _GEN_318 : _GEN_286; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_358 = _T_25 ? _GEN_319 : _GEN_287; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_359 = _T_25 ? _GEN_320 : _GEN_288; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_360 = _T_25 ? _GEN_321 : _GEN_289; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_361 = _T_25 ? _GEN_322 : _GEN_290; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_362 = _T_25 ? _GEN_323 : _GEN_291; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_363 = _T_25 ? _GEN_324 : _GEN_292; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_364 = _T_25 ? _GEN_325 : _GEN_293; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_365 = _T_25 ? _GEN_326 : _GEN_294; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_366 = _T_25 ? _GEN_327 : _GEN_295; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_367 = _T_25 ? _GEN_328 : _GEN_296; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_368 = _T_25 ? _GEN_329 : _GEN_297; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_369 = _T_25 ? _GEN_330 : _GEN_298; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_370 = _T_25 ? _GEN_331 : _GEN_299; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_371 = _T_25 ? _GEN_332 : _GEN_300; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_372 = _T_25 ? _GEN_333 : _GEN_301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_373 = _T_25 ? _GEN_334 : _GEN_302; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_374 = _T_25 ? _GEN_335 : _GEN_303; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_375 = _T_25 ? _GEN_336 : _GEN_304; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_376 = _T_25 ? _GEN_337 : _GEN_305; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_377 = _T_25 ? _GEN_338 : _GEN_306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_378 = _T_25 ? _GEN_339 : _GEN_307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_379 = _T_25 ? _GEN_340 : _GEN_308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_380 = _T_25 ? _GEN_341 : _GEN_309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_381 = _T_25 ? _GEN_342 : _GEN_310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_382 = _T_25 ? _GEN_343 : _GEN_311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_383 = _T_25 ? _GEN_344 : _GEN_312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_384 = _T_25 ? _GEN_345 : _GEN_313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_385 = _T_25 ? _GEN_346 : _GEN_314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_386 = _T_25 ? _GEN_347 : _GEN_315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _next_reg_T_10 = _GEN_31 ^ imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:62]
  wire [63:0] _GEN_388 = 5'h1 == rd ? _next_reg_T_10 : _GEN_356; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_389 = 5'h2 == rd ? _next_reg_T_10 : _GEN_357; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_390 = 5'h3 == rd ? _next_reg_T_10 : _GEN_358; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_391 = 5'h4 == rd ? _next_reg_T_10 : _GEN_359; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_392 = 5'h5 == rd ? _next_reg_T_10 : _GEN_360; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_393 = 5'h6 == rd ? _next_reg_T_10 : _GEN_361; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_394 = 5'h7 == rd ? _next_reg_T_10 : _GEN_362; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_395 = 5'h8 == rd ? _next_reg_T_10 : _GEN_363; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_396 = 5'h9 == rd ? _next_reg_T_10 : _GEN_364; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_397 = 5'ha == rd ? _next_reg_T_10 : _GEN_365; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_398 = 5'hb == rd ? _next_reg_T_10 : _GEN_366; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_399 = 5'hc == rd ? _next_reg_T_10 : _GEN_367; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_400 = 5'hd == rd ? _next_reg_T_10 : _GEN_368; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_401 = 5'he == rd ? _next_reg_T_10 : _GEN_369; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_402 = 5'hf == rd ? _next_reg_T_10 : _GEN_370; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_403 = 5'h10 == rd ? _next_reg_T_10 : _GEN_371; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_404 = 5'h11 == rd ? _next_reg_T_10 : _GEN_372; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_405 = 5'h12 == rd ? _next_reg_T_10 : _GEN_373; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_406 = 5'h13 == rd ? _next_reg_T_10 : _GEN_374; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_407 = 5'h14 == rd ? _next_reg_T_10 : _GEN_375; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_408 = 5'h15 == rd ? _next_reg_T_10 : _GEN_376; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_409 = 5'h16 == rd ? _next_reg_T_10 : _GEN_377; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_410 = 5'h17 == rd ? _next_reg_T_10 : _GEN_378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_411 = 5'h18 == rd ? _next_reg_T_10 : _GEN_379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_412 = 5'h19 == rd ? _next_reg_T_10 : _GEN_380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_413 = 5'h1a == rd ? _next_reg_T_10 : _GEN_381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_414 = 5'h1b == rd ? _next_reg_T_10 : _GEN_382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_415 = 5'h1c == rd ? _next_reg_T_10 : _GEN_383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_416 = 5'h1d == rd ? _next_reg_T_10 : _GEN_384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_417 = 5'h1e == rd ? _next_reg_T_10 : _GEN_385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_418 = 5'h1f == rd ? _next_reg_T_10 : _GEN_386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_427 = _T_31 ? _GEN_388 : _GEN_356; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_428 = _T_31 ? _GEN_389 : _GEN_357; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_429 = _T_31 ? _GEN_390 : _GEN_358; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_430 = _T_31 ? _GEN_391 : _GEN_359; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_431 = _T_31 ? _GEN_392 : _GEN_360; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_432 = _T_31 ? _GEN_393 : _GEN_361; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_433 = _T_31 ? _GEN_394 : _GEN_362; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_434 = _T_31 ? _GEN_395 : _GEN_363; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_435 = _T_31 ? _GEN_396 : _GEN_364; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_436 = _T_31 ? _GEN_397 : _GEN_365; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_437 = _T_31 ? _GEN_398 : _GEN_366; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_438 = _T_31 ? _GEN_399 : _GEN_367; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_439 = _T_31 ? _GEN_400 : _GEN_368; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_440 = _T_31 ? _GEN_401 : _GEN_369; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_441 = _T_31 ? _GEN_402 : _GEN_370; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_442 = _T_31 ? _GEN_403 : _GEN_371; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_443 = _T_31 ? _GEN_404 : _GEN_372; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_444 = _T_31 ? _GEN_405 : _GEN_373; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_445 = _T_31 ? _GEN_406 : _GEN_374; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_446 = _T_31 ? _GEN_407 : _GEN_375; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_447 = _T_31 ? _GEN_408 : _GEN_376; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_448 = _T_31 ? _GEN_409 : _GEN_377; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_449 = _T_31 ? _GEN_410 : _GEN_378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_450 = _T_31 ? _GEN_411 : _GEN_379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_451 = _T_31 ? _GEN_412 : _GEN_380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_452 = _T_31 ? _GEN_413 : _GEN_381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_453 = _T_31 ? _GEN_414 : _GEN_382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_454 = _T_31 ? _GEN_415 : _GEN_383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_455 = _T_31 ? _GEN_416 : _GEN_384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_456 = _T_31 ? _GEN_417 : _GEN_385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_457 = _T_31 ? _GEN_418 : _GEN_386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [94:0] _GEN_0 = {{31'd0}, _GEN_31}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:62]
  wire [94:0] _next_reg_T_12 = _GEN_0 << imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:62]
  wire [63:0] _GEN_459 = 5'h1 == rd ? _next_reg_T_12[63:0] : _GEN_427; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_460 = 5'h2 == rd ? _next_reg_T_12[63:0] : _GEN_428; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_461 = 5'h3 == rd ? _next_reg_T_12[63:0] : _GEN_429; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_462 = 5'h4 == rd ? _next_reg_T_12[63:0] : _GEN_430; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_463 = 5'h5 == rd ? _next_reg_T_12[63:0] : _GEN_431; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_464 = 5'h6 == rd ? _next_reg_T_12[63:0] : _GEN_432; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_465 = 5'h7 == rd ? _next_reg_T_12[63:0] : _GEN_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_466 = 5'h8 == rd ? _next_reg_T_12[63:0] : _GEN_434; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_467 = 5'h9 == rd ? _next_reg_T_12[63:0] : _GEN_435; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_468 = 5'ha == rd ? _next_reg_T_12[63:0] : _GEN_436; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_469 = 5'hb == rd ? _next_reg_T_12[63:0] : _GEN_437; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_470 = 5'hc == rd ? _next_reg_T_12[63:0] : _GEN_438; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_471 = 5'hd == rd ? _next_reg_T_12[63:0] : _GEN_439; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_472 = 5'he == rd ? _next_reg_T_12[63:0] : _GEN_440; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_473 = 5'hf == rd ? _next_reg_T_12[63:0] : _GEN_441; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_474 = 5'h10 == rd ? _next_reg_T_12[63:0] : _GEN_442; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_475 = 5'h11 == rd ? _next_reg_T_12[63:0] : _GEN_443; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_476 = 5'h12 == rd ? _next_reg_T_12[63:0] : _GEN_444; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_477 = 5'h13 == rd ? _next_reg_T_12[63:0] : _GEN_445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_478 = 5'h14 == rd ? _next_reg_T_12[63:0] : _GEN_446; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_479 = 5'h15 == rd ? _next_reg_T_12[63:0] : _GEN_447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_480 = 5'h16 == rd ? _next_reg_T_12[63:0] : _GEN_448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_481 = 5'h17 == rd ? _next_reg_T_12[63:0] : _GEN_449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_482 = 5'h18 == rd ? _next_reg_T_12[63:0] : _GEN_450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_483 = 5'h19 == rd ? _next_reg_T_12[63:0] : _GEN_451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_484 = 5'h1a == rd ? _next_reg_T_12[63:0] : _GEN_452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_485 = 5'h1b == rd ? _next_reg_T_12[63:0] : _GEN_453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_486 = 5'h1c == rd ? _next_reg_T_12[63:0] : _GEN_454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_487 = 5'h1d == rd ? _next_reg_T_12[63:0] : _GEN_455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_488 = 5'h1e == rd ? _next_reg_T_12[63:0] : _GEN_456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_489 = 5'h1f == rd ? _next_reg_T_12[63:0] : _GEN_457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_498 = _T_545 ? _GEN_459 : _GEN_427; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_499 = _T_545 ? _GEN_460 : _GEN_428; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_500 = _T_545 ? _GEN_461 : _GEN_429; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_501 = _T_545 ? _GEN_462 : _GEN_430; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_502 = _T_545 ? _GEN_463 : _GEN_431; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_503 = _T_545 ? _GEN_464 : _GEN_432; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_504 = _T_545 ? _GEN_465 : _GEN_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_505 = _T_545 ? _GEN_466 : _GEN_434; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_506 = _T_545 ? _GEN_467 : _GEN_435; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_507 = _T_545 ? _GEN_468 : _GEN_436; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_508 = _T_545 ? _GEN_469 : _GEN_437; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_509 = _T_545 ? _GEN_470 : _GEN_438; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_510 = _T_545 ? _GEN_471 : _GEN_439; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_511 = _T_545 ? _GEN_472 : _GEN_440; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_512 = _T_545 ? _GEN_473 : _GEN_441; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_513 = _T_545 ? _GEN_474 : _GEN_442; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_514 = _T_545 ? _GEN_475 : _GEN_443; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_515 = _T_545 ? _GEN_476 : _GEN_444; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_516 = _T_545 ? _GEN_477 : _GEN_445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_517 = _T_545 ? _GEN_478 : _GEN_446; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_518 = _T_545 ? _GEN_479 : _GEN_447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_519 = _T_545 ? _GEN_480 : _GEN_448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_520 = _T_545 ? _GEN_481 : _GEN_449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_521 = _T_545 ? _GEN_482 : _GEN_450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_522 = _T_545 ? _GEN_483 : _GEN_451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_523 = _T_545 ? _GEN_484 : _GEN_452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_524 = _T_545 ? _GEN_485 : _GEN_453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_525 = _T_545 ? _GEN_486 : _GEN_454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_526 = _T_545 ? _GEN_487 : _GEN_455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_527 = _T_545 ? _GEN_488 : _GEN_456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_528 = _T_545 ? _GEN_489 : _GEN_457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _next_reg_T_14 = _GEN_31 >> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:62]
  wire [63:0] _GEN_530 = 5'h1 == rd ? _next_reg_T_14 : _GEN_498; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_531 = 5'h2 == rd ? _next_reg_T_14 : _GEN_499; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_532 = 5'h3 == rd ? _next_reg_T_14 : _GEN_500; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_533 = 5'h4 == rd ? _next_reg_T_14 : _GEN_501; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_534 = 5'h5 == rd ? _next_reg_T_14 : _GEN_502; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_535 = 5'h6 == rd ? _next_reg_T_14 : _GEN_503; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_536 = 5'h7 == rd ? _next_reg_T_14 : _GEN_504; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_537 = 5'h8 == rd ? _next_reg_T_14 : _GEN_505; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_538 = 5'h9 == rd ? _next_reg_T_14 : _GEN_506; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_539 = 5'ha == rd ? _next_reg_T_14 : _GEN_507; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_540 = 5'hb == rd ? _next_reg_T_14 : _GEN_508; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_541 = 5'hc == rd ? _next_reg_T_14 : _GEN_509; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_542 = 5'hd == rd ? _next_reg_T_14 : _GEN_510; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_543 = 5'he == rd ? _next_reg_T_14 : _GEN_511; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_544 = 5'hf == rd ? _next_reg_T_14 : _GEN_512; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_545 = 5'h10 == rd ? _next_reg_T_14 : _GEN_513; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_546 = 5'h11 == rd ? _next_reg_T_14 : _GEN_514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_547 = 5'h12 == rd ? _next_reg_T_14 : _GEN_515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_548 = 5'h13 == rd ? _next_reg_T_14 : _GEN_516; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_549 = 5'h14 == rd ? _next_reg_T_14 : _GEN_517; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_550 = 5'h15 == rd ? _next_reg_T_14 : _GEN_518; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_551 = 5'h16 == rd ? _next_reg_T_14 : _GEN_519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_552 = 5'h17 == rd ? _next_reg_T_14 : _GEN_520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_553 = 5'h18 == rd ? _next_reg_T_14 : _GEN_521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_554 = 5'h19 == rd ? _next_reg_T_14 : _GEN_522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_555 = 5'h1a == rd ? _next_reg_T_14 : _GEN_523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_556 = 5'h1b == rd ? _next_reg_T_14 : _GEN_524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_557 = 5'h1c == rd ? _next_reg_T_14 : _GEN_525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_558 = 5'h1d == rd ? _next_reg_T_14 : _GEN_526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_559 = 5'h1e == rd ? _next_reg_T_14 : _GEN_527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_560 = 5'h1f == rd ? _next_reg_T_14 : _GEN_528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_569 = _T_551 ? _GEN_530 : _GEN_498; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_570 = _T_551 ? _GEN_531 : _GEN_499; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_571 = _T_551 ? _GEN_532 : _GEN_500; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_572 = _T_551 ? _GEN_533 : _GEN_501; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_573 = _T_551 ? _GEN_534 : _GEN_502; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_574 = _T_551 ? _GEN_535 : _GEN_503; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_575 = _T_551 ? _GEN_536 : _GEN_504; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_576 = _T_551 ? _GEN_537 : _GEN_505; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_577 = _T_551 ? _GEN_538 : _GEN_506; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_578 = _T_551 ? _GEN_539 : _GEN_507; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_579 = _T_551 ? _GEN_540 : _GEN_508; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_580 = _T_551 ? _GEN_541 : _GEN_509; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_581 = _T_551 ? _GEN_542 : _GEN_510; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_582 = _T_551 ? _GEN_543 : _GEN_511; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_583 = _T_551 ? _GEN_544 : _GEN_512; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_584 = _T_551 ? _GEN_545 : _GEN_513; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_585 = _T_551 ? _GEN_546 : _GEN_514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_586 = _T_551 ? _GEN_547 : _GEN_515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_587 = _T_551 ? _GEN_548 : _GEN_516; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_588 = _T_551 ? _GEN_549 : _GEN_517; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_589 = _T_551 ? _GEN_550 : _GEN_518; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_590 = _T_551 ? _GEN_551 : _GEN_519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_591 = _T_551 ? _GEN_552 : _GEN_520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_592 = _T_551 ? _GEN_553 : _GEN_521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_593 = _T_551 ? _GEN_554 : _GEN_522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_594 = _T_551 ? _GEN_555 : _GEN_523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_595 = _T_551 ? _GEN_556 : _GEN_524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_596 = _T_551 ? _GEN_557 : _GEN_525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_597 = _T_551 ? _GEN_558 : _GEN_526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_598 = _T_551 ? _GEN_559 : _GEN_527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_599 = _T_551 ? _GEN_560 : _GEN_528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _next_reg_T_18 = $signed(_T_300) >>> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:84]
  wire [63:0] _GEN_601 = 5'h1 == rd ? _next_reg_T_18 : _GEN_569; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_602 = 5'h2 == rd ? _next_reg_T_18 : _GEN_570; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_603 = 5'h3 == rd ? _next_reg_T_18 : _GEN_571; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_604 = 5'h4 == rd ? _next_reg_T_18 : _GEN_572; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_605 = 5'h5 == rd ? _next_reg_T_18 : _GEN_573; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_606 = 5'h6 == rd ? _next_reg_T_18 : _GEN_574; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_607 = 5'h7 == rd ? _next_reg_T_18 : _GEN_575; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_608 = 5'h8 == rd ? _next_reg_T_18 : _GEN_576; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_609 = 5'h9 == rd ? _next_reg_T_18 : _GEN_577; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_610 = 5'ha == rd ? _next_reg_T_18 : _GEN_578; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_611 = 5'hb == rd ? _next_reg_T_18 : _GEN_579; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_612 = 5'hc == rd ? _next_reg_T_18 : _GEN_580; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_613 = 5'hd == rd ? _next_reg_T_18 : _GEN_581; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_614 = 5'he == rd ? _next_reg_T_18 : _GEN_582; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_615 = 5'hf == rd ? _next_reg_T_18 : _GEN_583; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_616 = 5'h10 == rd ? _next_reg_T_18 : _GEN_584; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_617 = 5'h11 == rd ? _next_reg_T_18 : _GEN_585; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_618 = 5'h12 == rd ? _next_reg_T_18 : _GEN_586; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_619 = 5'h13 == rd ? _next_reg_T_18 : _GEN_587; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_620 = 5'h14 == rd ? _next_reg_T_18 : _GEN_588; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_621 = 5'h15 == rd ? _next_reg_T_18 : _GEN_589; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_622 = 5'h16 == rd ? _next_reg_T_18 : _GEN_590; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_623 = 5'h17 == rd ? _next_reg_T_18 : _GEN_591; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_624 = 5'h18 == rd ? _next_reg_T_18 : _GEN_592; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_625 = 5'h19 == rd ? _next_reg_T_18 : _GEN_593; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_626 = 5'h1a == rd ? _next_reg_T_18 : _GEN_594; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_627 = 5'h1b == rd ? _next_reg_T_18 : _GEN_595; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_628 = 5'h1c == rd ? _next_reg_T_18 : _GEN_596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_629 = 5'h1d == rd ? _next_reg_T_18 : _GEN_597; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_630 = 5'h1e == rd ? _next_reg_T_18 : _GEN_598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_631 = 5'h1f == rd ? _next_reg_T_18 : _GEN_599; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_640 = _T_557 ? _GEN_601 : _GEN_569; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_641 = _T_557 ? _GEN_602 : _GEN_570; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_642 = _T_557 ? _GEN_603 : _GEN_571; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_643 = _T_557 ? _GEN_604 : _GEN_572; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_644 = _T_557 ? _GEN_605 : _GEN_573; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_645 = _T_557 ? _GEN_606 : _GEN_574; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_646 = _T_557 ? _GEN_607 : _GEN_575; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_647 = _T_557 ? _GEN_608 : _GEN_576; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_648 = _T_557 ? _GEN_609 : _GEN_577; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_649 = _T_557 ? _GEN_610 : _GEN_578; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_650 = _T_557 ? _GEN_611 : _GEN_579; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_651 = _T_557 ? _GEN_612 : _GEN_580; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_652 = _T_557 ? _GEN_613 : _GEN_581; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_653 = _T_557 ? _GEN_614 : _GEN_582; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_654 = _T_557 ? _GEN_615 : _GEN_583; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_655 = _T_557 ? _GEN_616 : _GEN_584; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_656 = _T_557 ? _GEN_617 : _GEN_585; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_657 = _T_557 ? _GEN_618 : _GEN_586; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_658 = _T_557 ? _GEN_619 : _GEN_587; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_659 = _T_557 ? _GEN_620 : _GEN_588; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_660 = _T_557 ? _GEN_621 : _GEN_589; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_661 = _T_557 ? _GEN_622 : _GEN_590; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_662 = _T_557 ? _GEN_623 : _GEN_591; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_663 = _T_557 ? _GEN_624 : _GEN_592; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_664 = _T_557 ? _GEN_625 : _GEN_593; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_665 = _T_557 ? _GEN_626 : _GEN_594; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_666 = _T_557 ? _GEN_627 : _GEN_595; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_667 = _T_557 ? _GEN_628 : _GEN_596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_668 = _T_557 ? _GEN_629 : _GEN_597; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_669 = _T_557 ? _GEN_630 : _GEN_598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_670 = _T_557 ? _GEN_631 : _GEN_599; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_672 = 5'h1 == rd ? imm : _GEN_640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_673 = 5'h2 == rd ? imm : _GEN_641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_674 = 5'h3 == rd ? imm : _GEN_642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_675 = 5'h4 == rd ? imm : _GEN_643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_676 = 5'h5 == rd ? imm : _GEN_644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_677 = 5'h6 == rd ? imm : _GEN_645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_678 = 5'h7 == rd ? imm : _GEN_646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_679 = 5'h8 == rd ? imm : _GEN_647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_680 = 5'h9 == rd ? imm : _GEN_648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_681 = 5'ha == rd ? imm : _GEN_649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_682 = 5'hb == rd ? imm : _GEN_650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_683 = 5'hc == rd ? imm : _GEN_651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_684 = 5'hd == rd ? imm : _GEN_652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_685 = 5'he == rd ? imm : _GEN_653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_686 = 5'hf == rd ? imm : _GEN_654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_687 = 5'h10 == rd ? imm : _GEN_655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_688 = 5'h11 == rd ? imm : _GEN_656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_689 = 5'h12 == rd ? imm : _GEN_657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_690 = 5'h13 == rd ? imm : _GEN_658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_691 = 5'h14 == rd ? imm : _GEN_659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_692 = 5'h15 == rd ? imm : _GEN_660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_693 = 5'h16 == rd ? imm : _GEN_661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_694 = 5'h17 == rd ? imm : _GEN_662; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_695 = 5'h18 == rd ? imm : _GEN_663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_696 = 5'h19 == rd ? imm : _GEN_664; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_697 = 5'h1a == rd ? imm : _GEN_665; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_698 = 5'h1b == rd ? imm : _GEN_666; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_699 = 5'h1c == rd ? imm : _GEN_667; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_700 = 5'h1d == rd ? imm : _GEN_668; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_701 = 5'h1e == rd ? imm : _GEN_669; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_702 = 5'h1f == rd ? imm : _GEN_670; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_709 = _T_55 ? _GEN_672 : _GEN_640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_710 = _T_55 ? _GEN_673 : _GEN_641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_711 = _T_55 ? _GEN_674 : _GEN_642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_712 = _T_55 ? _GEN_675 : _GEN_643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_713 = _T_55 ? _GEN_676 : _GEN_644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_714 = _T_55 ? _GEN_677 : _GEN_645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_715 = _T_55 ? _GEN_678 : _GEN_646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_716 = _T_55 ? _GEN_679 : _GEN_647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_717 = _T_55 ? _GEN_680 : _GEN_648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_718 = _T_55 ? _GEN_681 : _GEN_649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_719 = _T_55 ? _GEN_682 : _GEN_650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_720 = _T_55 ? _GEN_683 : _GEN_651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_721 = _T_55 ? _GEN_684 : _GEN_652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_722 = _T_55 ? _GEN_685 : _GEN_653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_723 = _T_55 ? _GEN_686 : _GEN_654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_724 = _T_55 ? _GEN_687 : _GEN_655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_725 = _T_55 ? _GEN_688 : _GEN_656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_726 = _T_55 ? _GEN_689 : _GEN_657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_727 = _T_55 ? _GEN_690 : _GEN_658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_728 = _T_55 ? _GEN_691 : _GEN_659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_729 = _T_55 ? _GEN_692 : _GEN_660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_730 = _T_55 ? _GEN_693 : _GEN_661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_731 = _T_55 ? _GEN_694 : _GEN_662; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_732 = _T_55 ? _GEN_695 : _GEN_663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_733 = _T_55 ? _GEN_696 : _GEN_664; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_734 = _T_55 ? _GEN_697 : _GEN_665; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_735 = _T_55 ? _GEN_698 : _GEN_666; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_736 = _T_55 ? _GEN_699 : _GEN_667; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_737 = _T_55 ? _GEN_700 : _GEN_668; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_738 = _T_55 ? _GEN_701 : _GEN_669; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_739 = _T_55 ? _GEN_702 : _GEN_670; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_741 = 5'h1 == rd ? _T_334 : _GEN_709; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_742 = 5'h2 == rd ? _T_334 : _GEN_710; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_743 = 5'h3 == rd ? _T_334 : _GEN_711; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_744 = 5'h4 == rd ? _T_334 : _GEN_712; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_745 = 5'h5 == rd ? _T_334 : _GEN_713; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_746 = 5'h6 == rd ? _T_334 : _GEN_714; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_747 = 5'h7 == rd ? _T_334 : _GEN_715; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_748 = 5'h8 == rd ? _T_334 : _GEN_716; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_749 = 5'h9 == rd ? _T_334 : _GEN_717; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_750 = 5'ha == rd ? _T_334 : _GEN_718; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_751 = 5'hb == rd ? _T_334 : _GEN_719; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_752 = 5'hc == rd ? _T_334 : _GEN_720; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_753 = 5'hd == rd ? _T_334 : _GEN_721; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_754 = 5'he == rd ? _T_334 : _GEN_722; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_755 = 5'hf == rd ? _T_334 : _GEN_723; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_756 = 5'h10 == rd ? _T_334 : _GEN_724; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_757 = 5'h11 == rd ? _T_334 : _GEN_725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_758 = 5'h12 == rd ? _T_334 : _GEN_726; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_759 = 5'h13 == rd ? _T_334 : _GEN_727; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_760 = 5'h14 == rd ? _T_334 : _GEN_728; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_761 = 5'h15 == rd ? _T_334 : _GEN_729; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_762 = 5'h16 == rd ? _T_334 : _GEN_730; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_763 = 5'h17 == rd ? _T_334 : _GEN_731; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_764 = 5'h18 == rd ? _T_334 : _GEN_732; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_765 = 5'h19 == rd ? _T_334 : _GEN_733; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_766 = 5'h1a == rd ? _T_334 : _GEN_734; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_767 = 5'h1b == rd ? _T_334 : _GEN_735; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_768 = 5'h1c == rd ? _T_334 : _GEN_736; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_769 = 5'h1d == rd ? _T_334 : _GEN_737; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_770 = 5'h1e == rd ? _T_334 : _GEN_738; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_771 = 5'h1f == rd ? _T_334 : _GEN_739; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_778 = _T_59 ? _GEN_741 : _GEN_709; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_779 = _T_59 ? _GEN_742 : _GEN_710; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_780 = _T_59 ? _GEN_743 : _GEN_711; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_781 = _T_59 ? _GEN_744 : _GEN_712; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_782 = _T_59 ? _GEN_745 : _GEN_713; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_783 = _T_59 ? _GEN_746 : _GEN_714; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_784 = _T_59 ? _GEN_747 : _GEN_715; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_785 = _T_59 ? _GEN_748 : _GEN_716; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_786 = _T_59 ? _GEN_749 : _GEN_717; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_787 = _T_59 ? _GEN_750 : _GEN_718; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_788 = _T_59 ? _GEN_751 : _GEN_719; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_789 = _T_59 ? _GEN_752 : _GEN_720; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_790 = _T_59 ? _GEN_753 : _GEN_721; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_791 = _T_59 ? _GEN_754 : _GEN_722; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_792 = _T_59 ? _GEN_755 : _GEN_723; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_793 = _T_59 ? _GEN_756 : _GEN_724; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_794 = _T_59 ? _GEN_757 : _GEN_725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_795 = _T_59 ? _GEN_758 : _GEN_726; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_796 = _T_59 ? _GEN_759 : _GEN_727; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_797 = _T_59 ? _GEN_760 : _GEN_728; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_798 = _T_59 ? _GEN_761 : _GEN_729; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_799 = _T_59 ? _GEN_762 : _GEN_730; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_800 = _T_59 ? _GEN_763 : _GEN_731; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_801 = _T_59 ? _GEN_764 : _GEN_732; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_802 = _T_59 ? _GEN_765 : _GEN_733; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_803 = _T_59 ? _GEN_766 : _GEN_734; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_804 = _T_59 ? _GEN_767 : _GEN_735; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_805 = _T_59 ? _GEN_768 : _GEN_736; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_806 = _T_59 ? _GEN_769 : _GEN_737; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_807 = _T_59 ? _GEN_770 : _GEN_738; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_808 = _T_59 ? _GEN_771 : _GEN_739; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _next_reg_T_22 = _GEN_31 + _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:62]
  wire [63:0] _GEN_842 = 5'h1 == rd ? _next_reg_T_22 : _GEN_778; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_843 = 5'h2 == rd ? _next_reg_T_22 : _GEN_779; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_844 = 5'h3 == rd ? _next_reg_T_22 : _GEN_780; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_845 = 5'h4 == rd ? _next_reg_T_22 : _GEN_781; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_846 = 5'h5 == rd ? _next_reg_T_22 : _GEN_782; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_847 = 5'h6 == rd ? _next_reg_T_22 : _GEN_783; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_848 = 5'h7 == rd ? _next_reg_T_22 : _GEN_784; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_849 = 5'h8 == rd ? _next_reg_T_22 : _GEN_785; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_850 = 5'h9 == rd ? _next_reg_T_22 : _GEN_786; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_851 = 5'ha == rd ? _next_reg_T_22 : _GEN_787; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_852 = 5'hb == rd ? _next_reg_T_22 : _GEN_788; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_853 = 5'hc == rd ? _next_reg_T_22 : _GEN_789; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_854 = 5'hd == rd ? _next_reg_T_22 : _GEN_790; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_855 = 5'he == rd ? _next_reg_T_22 : _GEN_791; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_856 = 5'hf == rd ? _next_reg_T_22 : _GEN_792; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_857 = 5'h10 == rd ? _next_reg_T_22 : _GEN_793; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_858 = 5'h11 == rd ? _next_reg_T_22 : _GEN_794; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_859 = 5'h12 == rd ? _next_reg_T_22 : _GEN_795; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_860 = 5'h13 == rd ? _next_reg_T_22 : _GEN_796; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_861 = 5'h14 == rd ? _next_reg_T_22 : _GEN_797; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_862 = 5'h15 == rd ? _next_reg_T_22 : _GEN_798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_863 = 5'h16 == rd ? _next_reg_T_22 : _GEN_799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_864 = 5'h17 == rd ? _next_reg_T_22 : _GEN_800; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_865 = 5'h18 == rd ? _next_reg_T_22 : _GEN_801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_866 = 5'h19 == rd ? _next_reg_T_22 : _GEN_802; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_867 = 5'h1a == rd ? _next_reg_T_22 : _GEN_803; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_868 = 5'h1b == rd ? _next_reg_T_22 : _GEN_804; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_869 = 5'h1c == rd ? _next_reg_T_22 : _GEN_805; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_870 = 5'h1d == rd ? _next_reg_T_22 : _GEN_806; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_871 = 5'h1e == rd ? _next_reg_T_22 : _GEN_807; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_872 = 5'h1f == rd ? _next_reg_T_22 : _GEN_808; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_881 = _T_63 ? _GEN_842 : _GEN_778; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_882 = _T_63 ? _GEN_843 : _GEN_779; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_883 = _T_63 ? _GEN_844 : _GEN_780; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_884 = _T_63 ? _GEN_845 : _GEN_781; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_885 = _T_63 ? _GEN_846 : _GEN_782; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_886 = _T_63 ? _GEN_847 : _GEN_783; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_887 = _T_63 ? _GEN_848 : _GEN_784; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_888 = _T_63 ? _GEN_849 : _GEN_785; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_889 = _T_63 ? _GEN_850 : _GEN_786; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_890 = _T_63 ? _GEN_851 : _GEN_787; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_891 = _T_63 ? _GEN_852 : _GEN_788; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_892 = _T_63 ? _GEN_853 : _GEN_789; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_893 = _T_63 ? _GEN_854 : _GEN_790; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_894 = _T_63 ? _GEN_855 : _GEN_791; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_895 = _T_63 ? _GEN_856 : _GEN_792; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_896 = _T_63 ? _GEN_857 : _GEN_793; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_897 = _T_63 ? _GEN_858 : _GEN_794; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_898 = _T_63 ? _GEN_859 : _GEN_795; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_899 = _T_63 ? _GEN_860 : _GEN_796; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_900 = _T_63 ? _GEN_861 : _GEN_797; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_901 = _T_63 ? _GEN_862 : _GEN_798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_902 = _T_63 ? _GEN_863 : _GEN_799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_903 = _T_63 ? _GEN_864 : _GEN_800; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_904 = _T_63 ? _GEN_865 : _GEN_801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_905 = _T_63 ? _GEN_866 : _GEN_802; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_906 = _T_63 ? _GEN_867 : _GEN_803; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_907 = _T_63 ? _GEN_868 : _GEN_804; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_908 = _T_63 ? _GEN_869 : _GEN_805; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_909 = _T_63 ? _GEN_870 : _GEN_806; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_910 = _T_63 ? _GEN_871 : _GEN_807; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_911 = _T_63 ? _GEN_872 : _GEN_808; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _next_reg_rd_11 = {{63'd0}, _T_246}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_913 = 5'h1 == rd ? _next_reg_rd_11 : _GEN_881; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_914 = 5'h2 == rd ? _next_reg_rd_11 : _GEN_882; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_915 = 5'h3 == rd ? _next_reg_rd_11 : _GEN_883; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_916 = 5'h4 == rd ? _next_reg_rd_11 : _GEN_884; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_917 = 5'h5 == rd ? _next_reg_rd_11 : _GEN_885; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_918 = 5'h6 == rd ? _next_reg_rd_11 : _GEN_886; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_919 = 5'h7 == rd ? _next_reg_rd_11 : _GEN_887; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_920 = 5'h8 == rd ? _next_reg_rd_11 : _GEN_888; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_921 = 5'h9 == rd ? _next_reg_rd_11 : _GEN_889; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_922 = 5'ha == rd ? _next_reg_rd_11 : _GEN_890; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_923 = 5'hb == rd ? _next_reg_rd_11 : _GEN_891; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_924 = 5'hc == rd ? _next_reg_rd_11 : _GEN_892; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_925 = 5'hd == rd ? _next_reg_rd_11 : _GEN_893; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_926 = 5'he == rd ? _next_reg_rd_11 : _GEN_894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_927 = 5'hf == rd ? _next_reg_rd_11 : _GEN_895; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_928 = 5'h10 == rd ? _next_reg_rd_11 : _GEN_896; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_929 = 5'h11 == rd ? _next_reg_rd_11 : _GEN_897; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_930 = 5'h12 == rd ? _next_reg_rd_11 : _GEN_898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_931 = 5'h13 == rd ? _next_reg_rd_11 : _GEN_899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_932 = 5'h14 == rd ? _next_reg_rd_11 : _GEN_900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_933 = 5'h15 == rd ? _next_reg_rd_11 : _GEN_901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_934 = 5'h16 == rd ? _next_reg_rd_11 : _GEN_902; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_935 = 5'h17 == rd ? _next_reg_rd_11 : _GEN_903; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_936 = 5'h18 == rd ? _next_reg_rd_11 : _GEN_904; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_937 = 5'h19 == rd ? _next_reg_rd_11 : _GEN_905; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_938 = 5'h1a == rd ? _next_reg_rd_11 : _GEN_906; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_939 = 5'h1b == rd ? _next_reg_rd_11 : _GEN_907; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_940 = 5'h1c == rd ? _next_reg_rd_11 : _GEN_908; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_941 = 5'h1d == rd ? _next_reg_rd_11 : _GEN_909; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_942 = 5'h1e == rd ? _next_reg_rd_11 : _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_943 = 5'h1f == rd ? _next_reg_rd_11 : _GEN_911; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_952 = _T_70 ? _GEN_913 : _GEN_881; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_953 = _T_70 ? _GEN_914 : _GEN_882; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_954 = _T_70 ? _GEN_915 : _GEN_883; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_955 = _T_70 ? _GEN_916 : _GEN_884; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_956 = _T_70 ? _GEN_917 : _GEN_885; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_957 = _T_70 ? _GEN_918 : _GEN_886; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_958 = _T_70 ? _GEN_919 : _GEN_887; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_959 = _T_70 ? _GEN_920 : _GEN_888; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_960 = _T_70 ? _GEN_921 : _GEN_889; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_961 = _T_70 ? _GEN_922 : _GEN_890; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_962 = _T_70 ? _GEN_923 : _GEN_891; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_963 = _T_70 ? _GEN_924 : _GEN_892; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_964 = _T_70 ? _GEN_925 : _GEN_893; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_965 = _T_70 ? _GEN_926 : _GEN_894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_966 = _T_70 ? _GEN_927 : _GEN_895; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_967 = _T_70 ? _GEN_928 : _GEN_896; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_968 = _T_70 ? _GEN_929 : _GEN_897; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_969 = _T_70 ? _GEN_930 : _GEN_898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_970 = _T_70 ? _GEN_931 : _GEN_899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_971 = _T_70 ? _GEN_932 : _GEN_900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_972 = _T_70 ? _GEN_933 : _GEN_901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_973 = _T_70 ? _GEN_934 : _GEN_902; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_974 = _T_70 ? _GEN_935 : _GEN_903; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_975 = _T_70 ? _GEN_936 : _GEN_904; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_976 = _T_70 ? _GEN_937 : _GEN_905; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_977 = _T_70 ? _GEN_938 : _GEN_906; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_978 = _T_70 ? _GEN_939 : _GEN_907; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_979 = _T_70 ? _GEN_940 : _GEN_908; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_980 = _T_70 ? _GEN_941 : _GEN_909; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_981 = _T_70 ? _GEN_942 : _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_982 = _T_70 ? _GEN_943 : _GEN_911; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _next_reg_rd_12 = {{63'd0}, _T_273}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_984 = 5'h1 == rd ? _next_reg_rd_12 : _GEN_952; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_985 = 5'h2 == rd ? _next_reg_rd_12 : _GEN_953; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_986 = 5'h3 == rd ? _next_reg_rd_12 : _GEN_954; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_987 = 5'h4 == rd ? _next_reg_rd_12 : _GEN_955; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_988 = 5'h5 == rd ? _next_reg_rd_12 : _GEN_956; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_989 = 5'h6 == rd ? _next_reg_rd_12 : _GEN_957; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_990 = 5'h7 == rd ? _next_reg_rd_12 : _GEN_958; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_991 = 5'h8 == rd ? _next_reg_rd_12 : _GEN_959; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_992 = 5'h9 == rd ? _next_reg_rd_12 : _GEN_960; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_993 = 5'ha == rd ? _next_reg_rd_12 : _GEN_961; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_994 = 5'hb == rd ? _next_reg_rd_12 : _GEN_962; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_995 = 5'hc == rd ? _next_reg_rd_12 : _GEN_963; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_996 = 5'hd == rd ? _next_reg_rd_12 : _GEN_964; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_997 = 5'he == rd ? _next_reg_rd_12 : _GEN_965; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_998 = 5'hf == rd ? _next_reg_rd_12 : _GEN_966; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_999 = 5'h10 == rd ? _next_reg_rd_12 : _GEN_967; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1000 = 5'h11 == rd ? _next_reg_rd_12 : _GEN_968; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1001 = 5'h12 == rd ? _next_reg_rd_12 : _GEN_969; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1002 = 5'h13 == rd ? _next_reg_rd_12 : _GEN_970; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1003 = 5'h14 == rd ? _next_reg_rd_12 : _GEN_971; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1004 = 5'h15 == rd ? _next_reg_rd_12 : _GEN_972; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1005 = 5'h16 == rd ? _next_reg_rd_12 : _GEN_973; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1006 = 5'h17 == rd ? _next_reg_rd_12 : _GEN_974; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1007 = 5'h18 == rd ? _next_reg_rd_12 : _GEN_975; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1008 = 5'h19 == rd ? _next_reg_rd_12 : _GEN_976; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1009 = 5'h1a == rd ? _next_reg_rd_12 : _GEN_977; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1010 = 5'h1b == rd ? _next_reg_rd_12 : _GEN_978; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1011 = 5'h1c == rd ? _next_reg_rd_12 : _GEN_979; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1012 = 5'h1d == rd ? _next_reg_rd_12 : _GEN_980; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1013 = 5'h1e == rd ? _next_reg_rd_12 : _GEN_981; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1014 = 5'h1f == rd ? _next_reg_rd_12 : _GEN_982; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1023 = _T_77 ? _GEN_984 : _GEN_952; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1024 = _T_77 ? _GEN_985 : _GEN_953; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1025 = _T_77 ? _GEN_986 : _GEN_954; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1026 = _T_77 ? _GEN_987 : _GEN_955; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1027 = _T_77 ? _GEN_988 : _GEN_956; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1028 = _T_77 ? _GEN_989 : _GEN_957; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1029 = _T_77 ? _GEN_990 : _GEN_958; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1030 = _T_77 ? _GEN_991 : _GEN_959; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1031 = _T_77 ? _GEN_992 : _GEN_960; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1032 = _T_77 ? _GEN_993 : _GEN_961; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1033 = _T_77 ? _GEN_994 : _GEN_962; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1034 = _T_77 ? _GEN_995 : _GEN_963; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1035 = _T_77 ? _GEN_996 : _GEN_964; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1036 = _T_77 ? _GEN_997 : _GEN_965; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1037 = _T_77 ? _GEN_998 : _GEN_966; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1038 = _T_77 ? _GEN_999 : _GEN_967; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1039 = _T_77 ? _GEN_1000 : _GEN_968; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1040 = _T_77 ? _GEN_1001 : _GEN_969; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1041 = _T_77 ? _GEN_1002 : _GEN_970; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1042 = _T_77 ? _GEN_1003 : _GEN_971; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1043 = _T_77 ? _GEN_1004 : _GEN_972; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1044 = _T_77 ? _GEN_1005 : _GEN_973; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1045 = _T_77 ? _GEN_1006 : _GEN_974; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1046 = _T_77 ? _GEN_1007 : _GEN_975; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1047 = _T_77 ? _GEN_1008 : _GEN_976; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1048 = _T_77 ? _GEN_1009 : _GEN_977; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1049 = _T_77 ? _GEN_1010 : _GEN_978; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1050 = _T_77 ? _GEN_1011 : _GEN_979; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1051 = _T_77 ? _GEN_1012 : _GEN_980; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1052 = _T_77 ? _GEN_1013 : _GEN_981; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1053 = _T_77 ? _GEN_1014 : _GEN_982; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _next_reg_T_29 = _GEN_31 & _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:61]
  wire [63:0] _GEN_1055 = 5'h1 == rd ? _next_reg_T_29 : _GEN_1023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1056 = 5'h2 == rd ? _next_reg_T_29 : _GEN_1024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1057 = 5'h3 == rd ? _next_reg_T_29 : _GEN_1025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1058 = 5'h4 == rd ? _next_reg_T_29 : _GEN_1026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1059 = 5'h5 == rd ? _next_reg_T_29 : _GEN_1027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1060 = 5'h6 == rd ? _next_reg_T_29 : _GEN_1028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1061 = 5'h7 == rd ? _next_reg_T_29 : _GEN_1029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1062 = 5'h8 == rd ? _next_reg_T_29 : _GEN_1030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1063 = 5'h9 == rd ? _next_reg_T_29 : _GEN_1031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1064 = 5'ha == rd ? _next_reg_T_29 : _GEN_1032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1065 = 5'hb == rd ? _next_reg_T_29 : _GEN_1033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1066 = 5'hc == rd ? _next_reg_T_29 : _GEN_1034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1067 = 5'hd == rd ? _next_reg_T_29 : _GEN_1035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1068 = 5'he == rd ? _next_reg_T_29 : _GEN_1036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1069 = 5'hf == rd ? _next_reg_T_29 : _GEN_1037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1070 = 5'h10 == rd ? _next_reg_T_29 : _GEN_1038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1071 = 5'h11 == rd ? _next_reg_T_29 : _GEN_1039; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1072 = 5'h12 == rd ? _next_reg_T_29 : _GEN_1040; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1073 = 5'h13 == rd ? _next_reg_T_29 : _GEN_1041; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1074 = 5'h14 == rd ? _next_reg_T_29 : _GEN_1042; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1075 = 5'h15 == rd ? _next_reg_T_29 : _GEN_1043; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1076 = 5'h16 == rd ? _next_reg_T_29 : _GEN_1044; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1077 = 5'h17 == rd ? _next_reg_T_29 : _GEN_1045; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1078 = 5'h18 == rd ? _next_reg_T_29 : _GEN_1046; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1079 = 5'h19 == rd ? _next_reg_T_29 : _GEN_1047; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1080 = 5'h1a == rd ? _next_reg_T_29 : _GEN_1048; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1081 = 5'h1b == rd ? _next_reg_T_29 : _GEN_1049; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1082 = 5'h1c == rd ? _next_reg_T_29 : _GEN_1050; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1083 = 5'h1d == rd ? _next_reg_T_29 : _GEN_1051; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1084 = 5'h1e == rd ? _next_reg_T_29 : _GEN_1052; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1085 = 5'h1f == rd ? _next_reg_T_29 : _GEN_1053; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1094 = _T_84 ? _GEN_1055 : _GEN_1023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1095 = _T_84 ? _GEN_1056 : _GEN_1024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1096 = _T_84 ? _GEN_1057 : _GEN_1025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1097 = _T_84 ? _GEN_1058 : _GEN_1026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1098 = _T_84 ? _GEN_1059 : _GEN_1027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1099 = _T_84 ? _GEN_1060 : _GEN_1028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1100 = _T_84 ? _GEN_1061 : _GEN_1029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1101 = _T_84 ? _GEN_1062 : _GEN_1030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1102 = _T_84 ? _GEN_1063 : _GEN_1031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1103 = _T_84 ? _GEN_1064 : _GEN_1032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1104 = _T_84 ? _GEN_1065 : _GEN_1033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1105 = _T_84 ? _GEN_1066 : _GEN_1034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1106 = _T_84 ? _GEN_1067 : _GEN_1035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1107 = _T_84 ? _GEN_1068 : _GEN_1036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1108 = _T_84 ? _GEN_1069 : _GEN_1037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1109 = _T_84 ? _GEN_1070 : _GEN_1038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1110 = _T_84 ? _GEN_1071 : _GEN_1039; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1111 = _T_84 ? _GEN_1072 : _GEN_1040; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1112 = _T_84 ? _GEN_1073 : _GEN_1041; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1113 = _T_84 ? _GEN_1074 : _GEN_1042; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1114 = _T_84 ? _GEN_1075 : _GEN_1043; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1115 = _T_84 ? _GEN_1076 : _GEN_1044; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1116 = _T_84 ? _GEN_1077 : _GEN_1045; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1117 = _T_84 ? _GEN_1078 : _GEN_1046; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1118 = _T_84 ? _GEN_1079 : _GEN_1047; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1119 = _T_84 ? _GEN_1080 : _GEN_1048; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1120 = _T_84 ? _GEN_1081 : _GEN_1049; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1121 = _T_84 ? _GEN_1082 : _GEN_1050; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1122 = _T_84 ? _GEN_1083 : _GEN_1051; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1123 = _T_84 ? _GEN_1084 : _GEN_1052; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1124 = _T_84 ? _GEN_1085 : _GEN_1053; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _next_reg_T_30 = _GEN_31 | _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:61]
  wire [63:0] _GEN_1126 = 5'h1 == rd ? _next_reg_T_30 : _GEN_1094; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1127 = 5'h2 == rd ? _next_reg_T_30 : _GEN_1095; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1128 = 5'h3 == rd ? _next_reg_T_30 : _GEN_1096; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1129 = 5'h4 == rd ? _next_reg_T_30 : _GEN_1097; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1130 = 5'h5 == rd ? _next_reg_T_30 : _GEN_1098; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1131 = 5'h6 == rd ? _next_reg_T_30 : _GEN_1099; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1132 = 5'h7 == rd ? _next_reg_T_30 : _GEN_1100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1133 = 5'h8 == rd ? _next_reg_T_30 : _GEN_1101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1134 = 5'h9 == rd ? _next_reg_T_30 : _GEN_1102; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1135 = 5'ha == rd ? _next_reg_T_30 : _GEN_1103; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1136 = 5'hb == rd ? _next_reg_T_30 : _GEN_1104; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1137 = 5'hc == rd ? _next_reg_T_30 : _GEN_1105; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1138 = 5'hd == rd ? _next_reg_T_30 : _GEN_1106; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1139 = 5'he == rd ? _next_reg_T_30 : _GEN_1107; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1140 = 5'hf == rd ? _next_reg_T_30 : _GEN_1108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1141 = 5'h10 == rd ? _next_reg_T_30 : _GEN_1109; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1142 = 5'h11 == rd ? _next_reg_T_30 : _GEN_1110; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1143 = 5'h12 == rd ? _next_reg_T_30 : _GEN_1111; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1144 = 5'h13 == rd ? _next_reg_T_30 : _GEN_1112; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1145 = 5'h14 == rd ? _next_reg_T_30 : _GEN_1113; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1146 = 5'h15 == rd ? _next_reg_T_30 : _GEN_1114; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1147 = 5'h16 == rd ? _next_reg_T_30 : _GEN_1115; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1148 = 5'h17 == rd ? _next_reg_T_30 : _GEN_1116; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1149 = 5'h18 == rd ? _next_reg_T_30 : _GEN_1117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1150 = 5'h19 == rd ? _next_reg_T_30 : _GEN_1118; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1151 = 5'h1a == rd ? _next_reg_T_30 : _GEN_1119; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1152 = 5'h1b == rd ? _next_reg_T_30 : _GEN_1120; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1153 = 5'h1c == rd ? _next_reg_T_30 : _GEN_1121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1154 = 5'h1d == rd ? _next_reg_T_30 : _GEN_1122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1155 = 5'h1e == rd ? _next_reg_T_30 : _GEN_1123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1156 = 5'h1f == rd ? _next_reg_T_30 : _GEN_1124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1165 = _T_91 ? _GEN_1126 : _GEN_1094; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1166 = _T_91 ? _GEN_1127 : _GEN_1095; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1167 = _T_91 ? _GEN_1128 : _GEN_1096; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1168 = _T_91 ? _GEN_1129 : _GEN_1097; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1169 = _T_91 ? _GEN_1130 : _GEN_1098; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1170 = _T_91 ? _GEN_1131 : _GEN_1099; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1171 = _T_91 ? _GEN_1132 : _GEN_1100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1172 = _T_91 ? _GEN_1133 : _GEN_1101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1173 = _T_91 ? _GEN_1134 : _GEN_1102; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1174 = _T_91 ? _GEN_1135 : _GEN_1103; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1175 = _T_91 ? _GEN_1136 : _GEN_1104; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1176 = _T_91 ? _GEN_1137 : _GEN_1105; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1177 = _T_91 ? _GEN_1138 : _GEN_1106; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1178 = _T_91 ? _GEN_1139 : _GEN_1107; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1179 = _T_91 ? _GEN_1140 : _GEN_1108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1180 = _T_91 ? _GEN_1141 : _GEN_1109; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1181 = _T_91 ? _GEN_1142 : _GEN_1110; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1182 = _T_91 ? _GEN_1143 : _GEN_1111; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1183 = _T_91 ? _GEN_1144 : _GEN_1112; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1184 = _T_91 ? _GEN_1145 : _GEN_1113; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1185 = _T_91 ? _GEN_1146 : _GEN_1114; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1186 = _T_91 ? _GEN_1147 : _GEN_1115; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1187 = _T_91 ? _GEN_1148 : _GEN_1116; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1188 = _T_91 ? _GEN_1149 : _GEN_1117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1189 = _T_91 ? _GEN_1150 : _GEN_1118; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1190 = _T_91 ? _GEN_1151 : _GEN_1119; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1191 = _T_91 ? _GEN_1152 : _GEN_1120; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1192 = _T_91 ? _GEN_1153 : _GEN_1121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1193 = _T_91 ? _GEN_1154 : _GEN_1122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1194 = _T_91 ? _GEN_1155 : _GEN_1123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1195 = _T_91 ? _GEN_1156 : _GEN_1124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _next_reg_T_31 = _GEN_31 ^ _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:61]
  wire [63:0] _GEN_1197 = 5'h1 == rd ? _next_reg_T_31 : _GEN_1165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1198 = 5'h2 == rd ? _next_reg_T_31 : _GEN_1166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1199 = 5'h3 == rd ? _next_reg_T_31 : _GEN_1167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1200 = 5'h4 == rd ? _next_reg_T_31 : _GEN_1168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1201 = 5'h5 == rd ? _next_reg_T_31 : _GEN_1169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1202 = 5'h6 == rd ? _next_reg_T_31 : _GEN_1170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1203 = 5'h7 == rd ? _next_reg_T_31 : _GEN_1171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1204 = 5'h8 == rd ? _next_reg_T_31 : _GEN_1172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1205 = 5'h9 == rd ? _next_reg_T_31 : _GEN_1173; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1206 = 5'ha == rd ? _next_reg_T_31 : _GEN_1174; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1207 = 5'hb == rd ? _next_reg_T_31 : _GEN_1175; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1208 = 5'hc == rd ? _next_reg_T_31 : _GEN_1176; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1209 = 5'hd == rd ? _next_reg_T_31 : _GEN_1177; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1210 = 5'he == rd ? _next_reg_T_31 : _GEN_1178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1211 = 5'hf == rd ? _next_reg_T_31 : _GEN_1179; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1212 = 5'h10 == rd ? _next_reg_T_31 : _GEN_1180; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1213 = 5'h11 == rd ? _next_reg_T_31 : _GEN_1181; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1214 = 5'h12 == rd ? _next_reg_T_31 : _GEN_1182; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1215 = 5'h13 == rd ? _next_reg_T_31 : _GEN_1183; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1216 = 5'h14 == rd ? _next_reg_T_31 : _GEN_1184; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1217 = 5'h15 == rd ? _next_reg_T_31 : _GEN_1185; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1218 = 5'h16 == rd ? _next_reg_T_31 : _GEN_1186; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1219 = 5'h17 == rd ? _next_reg_T_31 : _GEN_1187; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1220 = 5'h18 == rd ? _next_reg_T_31 : _GEN_1188; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1221 = 5'h19 == rd ? _next_reg_T_31 : _GEN_1189; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1222 = 5'h1a == rd ? _next_reg_T_31 : _GEN_1190; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1223 = 5'h1b == rd ? _next_reg_T_31 : _GEN_1191; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1224 = 5'h1c == rd ? _next_reg_T_31 : _GEN_1192; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1225 = 5'h1d == rd ? _next_reg_T_31 : _GEN_1193; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1226 = 5'h1e == rd ? _next_reg_T_31 : _GEN_1194; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1227 = 5'h1f == rd ? _next_reg_T_31 : _GEN_1195; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1236 = _T_98 ? _GEN_1197 : _GEN_1165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1237 = _T_98 ? _GEN_1198 : _GEN_1166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1238 = _T_98 ? _GEN_1199 : _GEN_1167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1239 = _T_98 ? _GEN_1200 : _GEN_1168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1240 = _T_98 ? _GEN_1201 : _GEN_1169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1241 = _T_98 ? _GEN_1202 : _GEN_1170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1242 = _T_98 ? _GEN_1203 : _GEN_1171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1243 = _T_98 ? _GEN_1204 : _GEN_1172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1244 = _T_98 ? _GEN_1205 : _GEN_1173; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1245 = _T_98 ? _GEN_1206 : _GEN_1174; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1246 = _T_98 ? _GEN_1207 : _GEN_1175; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1247 = _T_98 ? _GEN_1208 : _GEN_1176; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1248 = _T_98 ? _GEN_1209 : _GEN_1177; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1249 = _T_98 ? _GEN_1210 : _GEN_1178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1250 = _T_98 ? _GEN_1211 : _GEN_1179; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1251 = _T_98 ? _GEN_1212 : _GEN_1180; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1252 = _T_98 ? _GEN_1213 : _GEN_1181; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1253 = _T_98 ? _GEN_1214 : _GEN_1182; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1254 = _T_98 ? _GEN_1215 : _GEN_1183; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1255 = _T_98 ? _GEN_1216 : _GEN_1184; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1256 = _T_98 ? _GEN_1217 : _GEN_1185; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1257 = _T_98 ? _GEN_1218 : _GEN_1186; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1258 = _T_98 ? _GEN_1219 : _GEN_1187; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1259 = _T_98 ? _GEN_1220 : _GEN_1188; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1260 = _T_98 ? _GEN_1221 : _GEN_1189; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1261 = _T_98 ? _GEN_1222 : _GEN_1190; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1262 = _T_98 ? _GEN_1223 : _GEN_1191; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1263 = _T_98 ? _GEN_1224 : _GEN_1192; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1264 = _T_98 ? _GEN_1225 : _GEN_1193; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1265 = _T_98 ? _GEN_1226 : _GEN_1194; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1266 = _T_98 ? _GEN_1227 : _GEN_1195; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [94:0] _GEN_32 = {{31'd0}, _GEN_31}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:61]
  wire [94:0] _next_reg_T_33 = _GEN_32 << _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:61]
  wire [63:0] _GEN_1268 = 5'h1 == rd ? _next_reg_T_33[63:0] : _GEN_1236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1269 = 5'h2 == rd ? _next_reg_T_33[63:0] : _GEN_1237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1270 = 5'h3 == rd ? _next_reg_T_33[63:0] : _GEN_1238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1271 = 5'h4 == rd ? _next_reg_T_33[63:0] : _GEN_1239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1272 = 5'h5 == rd ? _next_reg_T_33[63:0] : _GEN_1240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1273 = 5'h6 == rd ? _next_reg_T_33[63:0] : _GEN_1241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1274 = 5'h7 == rd ? _next_reg_T_33[63:0] : _GEN_1242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1275 = 5'h8 == rd ? _next_reg_T_33[63:0] : _GEN_1243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1276 = 5'h9 == rd ? _next_reg_T_33[63:0] : _GEN_1244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1277 = 5'ha == rd ? _next_reg_T_33[63:0] : _GEN_1245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1278 = 5'hb == rd ? _next_reg_T_33[63:0] : _GEN_1246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1279 = 5'hc == rd ? _next_reg_T_33[63:0] : _GEN_1247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1280 = 5'hd == rd ? _next_reg_T_33[63:0] : _GEN_1248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1281 = 5'he == rd ? _next_reg_T_33[63:0] : _GEN_1249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1282 = 5'hf == rd ? _next_reg_T_33[63:0] : _GEN_1250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1283 = 5'h10 == rd ? _next_reg_T_33[63:0] : _GEN_1251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1284 = 5'h11 == rd ? _next_reg_T_33[63:0] : _GEN_1252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1285 = 5'h12 == rd ? _next_reg_T_33[63:0] : _GEN_1253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1286 = 5'h13 == rd ? _next_reg_T_33[63:0] : _GEN_1254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1287 = 5'h14 == rd ? _next_reg_T_33[63:0] : _GEN_1255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1288 = 5'h15 == rd ? _next_reg_T_33[63:0] : _GEN_1256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1289 = 5'h16 == rd ? _next_reg_T_33[63:0] : _GEN_1257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1290 = 5'h17 == rd ? _next_reg_T_33[63:0] : _GEN_1258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1291 = 5'h18 == rd ? _next_reg_T_33[63:0] : _GEN_1259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1292 = 5'h19 == rd ? _next_reg_T_33[63:0] : _GEN_1260; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1293 = 5'h1a == rd ? _next_reg_T_33[63:0] : _GEN_1261; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1294 = 5'h1b == rd ? _next_reg_T_33[63:0] : _GEN_1262; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1295 = 5'h1c == rd ? _next_reg_T_33[63:0] : _GEN_1263; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1296 = 5'h1d == rd ? _next_reg_T_33[63:0] : _GEN_1264; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1297 = 5'h1e == rd ? _next_reg_T_33[63:0] : _GEN_1265; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1298 = 5'h1f == rd ? _next_reg_T_33[63:0] : _GEN_1266; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1307 = _T_581 ? _GEN_1268 : _GEN_1236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1308 = _T_581 ? _GEN_1269 : _GEN_1237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1309 = _T_581 ? _GEN_1270 : _GEN_1238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1310 = _T_581 ? _GEN_1271 : _GEN_1239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1311 = _T_581 ? _GEN_1272 : _GEN_1240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1312 = _T_581 ? _GEN_1273 : _GEN_1241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1313 = _T_581 ? _GEN_1274 : _GEN_1242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1314 = _T_581 ? _GEN_1275 : _GEN_1243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1315 = _T_581 ? _GEN_1276 : _GEN_1244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1316 = _T_581 ? _GEN_1277 : _GEN_1245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1317 = _T_581 ? _GEN_1278 : _GEN_1246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1318 = _T_581 ? _GEN_1279 : _GEN_1247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1319 = _T_581 ? _GEN_1280 : _GEN_1248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1320 = _T_581 ? _GEN_1281 : _GEN_1249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1321 = _T_581 ? _GEN_1282 : _GEN_1250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1322 = _T_581 ? _GEN_1283 : _GEN_1251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1323 = _T_581 ? _GEN_1284 : _GEN_1252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1324 = _T_581 ? _GEN_1285 : _GEN_1253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1325 = _T_581 ? _GEN_1286 : _GEN_1254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1326 = _T_581 ? _GEN_1287 : _GEN_1255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1327 = _T_581 ? _GEN_1288 : _GEN_1256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1328 = _T_581 ? _GEN_1289 : _GEN_1257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1329 = _T_581 ? _GEN_1290 : _GEN_1258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1330 = _T_581 ? _GEN_1291 : _GEN_1259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1331 = _T_581 ? _GEN_1292 : _GEN_1260; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1332 = _T_581 ? _GEN_1293 : _GEN_1261; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1333 = _T_581 ? _GEN_1294 : _GEN_1262; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1334 = _T_581 ? _GEN_1295 : _GEN_1263; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1335 = _T_581 ? _GEN_1296 : _GEN_1264; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1336 = _T_581 ? _GEN_1297 : _GEN_1265; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1337 = _T_581 ? _GEN_1298 : _GEN_1266; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _next_reg_T_35 = _GEN_31 >> _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:61]
  wire [63:0] _GEN_1339 = 5'h1 == rd ? _next_reg_T_35 : _GEN_1307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1340 = 5'h2 == rd ? _next_reg_T_35 : _GEN_1308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1341 = 5'h3 == rd ? _next_reg_T_35 : _GEN_1309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1342 = 5'h4 == rd ? _next_reg_T_35 : _GEN_1310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1343 = 5'h5 == rd ? _next_reg_T_35 : _GEN_1311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1344 = 5'h6 == rd ? _next_reg_T_35 : _GEN_1312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1345 = 5'h7 == rd ? _next_reg_T_35 : _GEN_1313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1346 = 5'h8 == rd ? _next_reg_T_35 : _GEN_1314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1347 = 5'h9 == rd ? _next_reg_T_35 : _GEN_1315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1348 = 5'ha == rd ? _next_reg_T_35 : _GEN_1316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1349 = 5'hb == rd ? _next_reg_T_35 : _GEN_1317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1350 = 5'hc == rd ? _next_reg_T_35 : _GEN_1318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1351 = 5'hd == rd ? _next_reg_T_35 : _GEN_1319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1352 = 5'he == rd ? _next_reg_T_35 : _GEN_1320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1353 = 5'hf == rd ? _next_reg_T_35 : _GEN_1321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1354 = 5'h10 == rd ? _next_reg_T_35 : _GEN_1322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1355 = 5'h11 == rd ? _next_reg_T_35 : _GEN_1323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1356 = 5'h12 == rd ? _next_reg_T_35 : _GEN_1324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1357 = 5'h13 == rd ? _next_reg_T_35 : _GEN_1325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1358 = 5'h14 == rd ? _next_reg_T_35 : _GEN_1326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1359 = 5'h15 == rd ? _next_reg_T_35 : _GEN_1327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1360 = 5'h16 == rd ? _next_reg_T_35 : _GEN_1328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1361 = 5'h17 == rd ? _next_reg_T_35 : _GEN_1329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1362 = 5'h18 == rd ? _next_reg_T_35 : _GEN_1330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1363 = 5'h19 == rd ? _next_reg_T_35 : _GEN_1331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1364 = 5'h1a == rd ? _next_reg_T_35 : _GEN_1332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1365 = 5'h1b == rd ? _next_reg_T_35 : _GEN_1333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1366 = 5'h1c == rd ? _next_reg_T_35 : _GEN_1334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1367 = 5'h1d == rd ? _next_reg_T_35 : _GEN_1335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1368 = 5'h1e == rd ? _next_reg_T_35 : _GEN_1336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1369 = 5'h1f == rd ? _next_reg_T_35 : _GEN_1337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1378 = _T_588 ? _GEN_1339 : _GEN_1307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1379 = _T_588 ? _GEN_1340 : _GEN_1308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1380 = _T_588 ? _GEN_1341 : _GEN_1309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1381 = _T_588 ? _GEN_1342 : _GEN_1310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1382 = _T_588 ? _GEN_1343 : _GEN_1311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1383 = _T_588 ? _GEN_1344 : _GEN_1312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1384 = _T_588 ? _GEN_1345 : _GEN_1313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1385 = _T_588 ? _GEN_1346 : _GEN_1314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1386 = _T_588 ? _GEN_1347 : _GEN_1315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1387 = _T_588 ? _GEN_1348 : _GEN_1316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1388 = _T_588 ? _GEN_1349 : _GEN_1317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1389 = _T_588 ? _GEN_1350 : _GEN_1318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1390 = _T_588 ? _GEN_1351 : _GEN_1319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1391 = _T_588 ? _GEN_1352 : _GEN_1320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1392 = _T_588 ? _GEN_1353 : _GEN_1321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1393 = _T_588 ? _GEN_1354 : _GEN_1322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1394 = _T_588 ? _GEN_1355 : _GEN_1323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1395 = _T_588 ? _GEN_1356 : _GEN_1324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1396 = _T_588 ? _GEN_1357 : _GEN_1325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1397 = _T_588 ? _GEN_1358 : _GEN_1326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1398 = _T_588 ? _GEN_1359 : _GEN_1327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1399 = _T_588 ? _GEN_1360 : _GEN_1328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1400 = _T_588 ? _GEN_1361 : _GEN_1329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1401 = _T_588 ? _GEN_1362 : _GEN_1330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1402 = _T_588 ? _GEN_1363 : _GEN_1331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1403 = _T_588 ? _GEN_1364 : _GEN_1332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1404 = _T_588 ? _GEN_1365 : _GEN_1333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1405 = _T_588 ? _GEN_1366 : _GEN_1334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1406 = _T_588 ? _GEN_1367 : _GEN_1335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1407 = _T_588 ? _GEN_1368 : _GEN_1336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1408 = _T_588 ? _GEN_1369 : _GEN_1337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _next_reg_T_37 = _GEN_31 - _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:61]
  wire [63:0] _GEN_1410 = 5'h1 == rd ? _next_reg_T_37 : _GEN_1378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1411 = 5'h2 == rd ? _next_reg_T_37 : _GEN_1379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1412 = 5'h3 == rd ? _next_reg_T_37 : _GEN_1380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1413 = 5'h4 == rd ? _next_reg_T_37 : _GEN_1381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1414 = 5'h5 == rd ? _next_reg_T_37 : _GEN_1382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1415 = 5'h6 == rd ? _next_reg_T_37 : _GEN_1383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1416 = 5'h7 == rd ? _next_reg_T_37 : _GEN_1384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1417 = 5'h8 == rd ? _next_reg_T_37 : _GEN_1385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1418 = 5'h9 == rd ? _next_reg_T_37 : _GEN_1386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1419 = 5'ha == rd ? _next_reg_T_37 : _GEN_1387; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1420 = 5'hb == rd ? _next_reg_T_37 : _GEN_1388; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1421 = 5'hc == rd ? _next_reg_T_37 : _GEN_1389; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1422 = 5'hd == rd ? _next_reg_T_37 : _GEN_1390; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1423 = 5'he == rd ? _next_reg_T_37 : _GEN_1391; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1424 = 5'hf == rd ? _next_reg_T_37 : _GEN_1392; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1425 = 5'h10 == rd ? _next_reg_T_37 : _GEN_1393; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1426 = 5'h11 == rd ? _next_reg_T_37 : _GEN_1394; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1427 = 5'h12 == rd ? _next_reg_T_37 : _GEN_1395; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1428 = 5'h13 == rd ? _next_reg_T_37 : _GEN_1396; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1429 = 5'h14 == rd ? _next_reg_T_37 : _GEN_1397; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1430 = 5'h15 == rd ? _next_reg_T_37 : _GEN_1398; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1431 = 5'h16 == rd ? _next_reg_T_37 : _GEN_1399; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1432 = 5'h17 == rd ? _next_reg_T_37 : _GEN_1400; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1433 = 5'h18 == rd ? _next_reg_T_37 : _GEN_1401; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1434 = 5'h19 == rd ? _next_reg_T_37 : _GEN_1402; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1435 = 5'h1a == rd ? _next_reg_T_37 : _GEN_1403; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1436 = 5'h1b == rd ? _next_reg_T_37 : _GEN_1404; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1437 = 5'h1c == rd ? _next_reg_T_37 : _GEN_1405; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1438 = 5'h1d == rd ? _next_reg_T_37 : _GEN_1406; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1439 = 5'h1e == rd ? _next_reg_T_37 : _GEN_1407; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1440 = 5'h1f == rd ? _next_reg_T_37 : _GEN_1408; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1449 = _T_119 ? _GEN_1410 : _GEN_1378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1450 = _T_119 ? _GEN_1411 : _GEN_1379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1451 = _T_119 ? _GEN_1412 : _GEN_1380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1452 = _T_119 ? _GEN_1413 : _GEN_1381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1453 = _T_119 ? _GEN_1414 : _GEN_1382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1454 = _T_119 ? _GEN_1415 : _GEN_1383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1455 = _T_119 ? _GEN_1416 : _GEN_1384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1456 = _T_119 ? _GEN_1417 : _GEN_1385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1457 = _T_119 ? _GEN_1418 : _GEN_1386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1458 = _T_119 ? _GEN_1419 : _GEN_1387; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1459 = _T_119 ? _GEN_1420 : _GEN_1388; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1460 = _T_119 ? _GEN_1421 : _GEN_1389; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1461 = _T_119 ? _GEN_1422 : _GEN_1390; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1462 = _T_119 ? _GEN_1423 : _GEN_1391; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1463 = _T_119 ? _GEN_1424 : _GEN_1392; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1464 = _T_119 ? _GEN_1425 : _GEN_1393; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1465 = _T_119 ? _GEN_1426 : _GEN_1394; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1466 = _T_119 ? _GEN_1427 : _GEN_1395; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1467 = _T_119 ? _GEN_1428 : _GEN_1396; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1468 = _T_119 ? _GEN_1429 : _GEN_1397; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1469 = _T_119 ? _GEN_1430 : _GEN_1398; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1470 = _T_119 ? _GEN_1431 : _GEN_1399; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1471 = _T_119 ? _GEN_1432 : _GEN_1400; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1472 = _T_119 ? _GEN_1433 : _GEN_1401; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1473 = _T_119 ? _GEN_1434 : _GEN_1402; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1474 = _T_119 ? _GEN_1435 : _GEN_1403; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1475 = _T_119 ? _GEN_1436 : _GEN_1404; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1476 = _T_119 ? _GEN_1437 : _GEN_1405; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1477 = _T_119 ? _GEN_1438 : _GEN_1406; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1478 = _T_119 ? _GEN_1439 : _GEN_1407; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1479 = _T_119 ? _GEN_1440 : _GEN_1408; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _next_reg_T_41 = $signed(_T_300) >>> _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:92]
  wire [63:0] _GEN_1481 = 5'h1 == rd ? _next_reg_T_41 : _GEN_1449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1482 = 5'h2 == rd ? _next_reg_T_41 : _GEN_1450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1483 = 5'h3 == rd ? _next_reg_T_41 : _GEN_1451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1484 = 5'h4 == rd ? _next_reg_T_41 : _GEN_1452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1485 = 5'h5 == rd ? _next_reg_T_41 : _GEN_1453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1486 = 5'h6 == rd ? _next_reg_T_41 : _GEN_1454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1487 = 5'h7 == rd ? _next_reg_T_41 : _GEN_1455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1488 = 5'h8 == rd ? _next_reg_T_41 : _GEN_1456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1489 = 5'h9 == rd ? _next_reg_T_41 : _GEN_1457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1490 = 5'ha == rd ? _next_reg_T_41 : _GEN_1458; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1491 = 5'hb == rd ? _next_reg_T_41 : _GEN_1459; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1492 = 5'hc == rd ? _next_reg_T_41 : _GEN_1460; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1493 = 5'hd == rd ? _next_reg_T_41 : _GEN_1461; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1494 = 5'he == rd ? _next_reg_T_41 : _GEN_1462; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1495 = 5'hf == rd ? _next_reg_T_41 : _GEN_1463; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1496 = 5'h10 == rd ? _next_reg_T_41 : _GEN_1464; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1497 = 5'h11 == rd ? _next_reg_T_41 : _GEN_1465; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1498 = 5'h12 == rd ? _next_reg_T_41 : _GEN_1466; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1499 = 5'h13 == rd ? _next_reg_T_41 : _GEN_1467; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1500 = 5'h14 == rd ? _next_reg_T_41 : _GEN_1468; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1501 = 5'h15 == rd ? _next_reg_T_41 : _GEN_1469; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1502 = 5'h16 == rd ? _next_reg_T_41 : _GEN_1470; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1503 = 5'h17 == rd ? _next_reg_T_41 : _GEN_1471; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1504 = 5'h18 == rd ? _next_reg_T_41 : _GEN_1472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1505 = 5'h19 == rd ? _next_reg_T_41 : _GEN_1473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1506 = 5'h1a == rd ? _next_reg_T_41 : _GEN_1474; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1507 = 5'h1b == rd ? _next_reg_T_41 : _GEN_1475; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1508 = 5'h1c == rd ? _next_reg_T_41 : _GEN_1476; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1509 = 5'h1d == rd ? _next_reg_T_41 : _GEN_1477; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1510 = 5'h1e == rd ? _next_reg_T_41 : _GEN_1478; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1511 = 5'h1f == rd ? _next_reg_T_41 : _GEN_1479; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1520 = _T_595 ? _GEN_1481 : _GEN_1449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1521 = _T_595 ? _GEN_1482 : _GEN_1450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1522 = _T_595 ? _GEN_1483 : _GEN_1451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1523 = _T_595 ? _GEN_1484 : _GEN_1452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1524 = _T_595 ? _GEN_1485 : _GEN_1453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1525 = _T_595 ? _GEN_1486 : _GEN_1454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1526 = _T_595 ? _GEN_1487 : _GEN_1455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1527 = _T_595 ? _GEN_1488 : _GEN_1456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1528 = _T_595 ? _GEN_1489 : _GEN_1457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1529 = _T_595 ? _GEN_1490 : _GEN_1458; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1530 = _T_595 ? _GEN_1491 : _GEN_1459; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1531 = _T_595 ? _GEN_1492 : _GEN_1460; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1532 = _T_595 ? _GEN_1493 : _GEN_1461; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1533 = _T_595 ? _GEN_1494 : _GEN_1462; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1534 = _T_595 ? _GEN_1495 : _GEN_1463; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1535 = _T_595 ? _GEN_1496 : _GEN_1464; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1536 = _T_595 ? _GEN_1497 : _GEN_1465; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1537 = _T_595 ? _GEN_1498 : _GEN_1466; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1538 = _T_595 ? _GEN_1499 : _GEN_1467; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1539 = _T_595 ? _GEN_1500 : _GEN_1468; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1540 = _T_595 ? _GEN_1501 : _GEN_1469; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1541 = _T_595 ? _GEN_1502 : _GEN_1470; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1542 = _T_595 ? _GEN_1503 : _GEN_1471; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1543 = _T_595 ? _GEN_1504 : _GEN_1472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1544 = _T_595 ? _GEN_1505 : _GEN_1473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1545 = _T_595 ? _GEN_1506 : _GEN_1474; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1546 = _T_595 ? _GEN_1507 : _GEN_1475; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1547 = _T_595 ? _GEN_1508 : _GEN_1476; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1548 = _T_595 ? _GEN_1509 : _GEN_1477; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1549 = _T_595 ? _GEN_1510 : _GEN_1478; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1550 = _T_595 ? _GEN_1511 : _GEN_1479; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _next_reg_T_43 = io_now_pc + 64'h4; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:37]
  wire [63:0] _GEN_1552 = 5'h1 == rd ? _next_reg_T_43 : _GEN_1520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1553 = 5'h2 == rd ? _next_reg_T_43 : _GEN_1521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1554 = 5'h3 == rd ? _next_reg_T_43 : _GEN_1522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1555 = 5'h4 == rd ? _next_reg_T_43 : _GEN_1523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1556 = 5'h5 == rd ? _next_reg_T_43 : _GEN_1524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1557 = 5'h6 == rd ? _next_reg_T_43 : _GEN_1525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1558 = 5'h7 == rd ? _next_reg_T_43 : _GEN_1526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1559 = 5'h8 == rd ? _next_reg_T_43 : _GEN_1527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1560 = 5'h9 == rd ? _next_reg_T_43 : _GEN_1528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1561 = 5'ha == rd ? _next_reg_T_43 : _GEN_1529; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1562 = 5'hb == rd ? _next_reg_T_43 : _GEN_1530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1563 = 5'hc == rd ? _next_reg_T_43 : _GEN_1531; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1564 = 5'hd == rd ? _next_reg_T_43 : _GEN_1532; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1565 = 5'he == rd ? _next_reg_T_43 : _GEN_1533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1566 = 5'hf == rd ? _next_reg_T_43 : _GEN_1534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1567 = 5'h10 == rd ? _next_reg_T_43 : _GEN_1535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1568 = 5'h11 == rd ? _next_reg_T_43 : _GEN_1536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1569 = 5'h12 == rd ? _next_reg_T_43 : _GEN_1537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1570 = 5'h13 == rd ? _next_reg_T_43 : _GEN_1538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1571 = 5'h14 == rd ? _next_reg_T_43 : _GEN_1539; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1572 = 5'h15 == rd ? _next_reg_T_43 : _GEN_1540; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1573 = 5'h16 == rd ? _next_reg_T_43 : _GEN_1541; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1574 = 5'h17 == rd ? _next_reg_T_43 : _GEN_1542; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1575 = 5'h18 == rd ? _next_reg_T_43 : _GEN_1543; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1576 = 5'h19 == rd ? _next_reg_T_43 : _GEN_1544; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1577 = 5'h1a == rd ? _next_reg_T_43 : _GEN_1545; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1578 = 5'h1b == rd ? _next_reg_T_43 : _GEN_1546; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1579 = 5'h1c == rd ? _next_reg_T_43 : _GEN_1547; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1580 = 5'h1d == rd ? _next_reg_T_43 : _GEN_1548; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1581 = 5'h1e == rd ? _next_reg_T_43 : _GEN_1549; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1582 = 5'h1f == rd ? _next_reg_T_43 : _GEN_1550; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1584 = _T_346 ? _T_334 : io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55 191:27]
  wire [63:0] _GEN_1586 = _T_346 ? _GEN_1552 : _GEN_1520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1587 = _T_346 ? _GEN_1553 : _GEN_1521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1588 = _T_346 ? _GEN_1554 : _GEN_1522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1589 = _T_346 ? _GEN_1555 : _GEN_1523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1590 = _T_346 ? _GEN_1556 : _GEN_1524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1591 = _T_346 ? _GEN_1557 : _GEN_1525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1592 = _T_346 ? _GEN_1558 : _GEN_1526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1593 = _T_346 ? _GEN_1559 : _GEN_1527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1594 = _T_346 ? _GEN_1560 : _GEN_1528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1595 = _T_346 ? _GEN_1561 : _GEN_1529; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1596 = _T_346 ? _GEN_1562 : _GEN_1530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1597 = _T_346 ? _GEN_1563 : _GEN_1531; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1598 = _T_346 ? _GEN_1564 : _GEN_1532; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1599 = _T_346 ? _GEN_1565 : _GEN_1533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1600 = _T_346 ? _GEN_1566 : _GEN_1534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1601 = _T_346 ? _GEN_1567 : _GEN_1535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1602 = _T_346 ? _GEN_1568 : _GEN_1536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1603 = _T_346 ? _GEN_1569 : _GEN_1537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1604 = _T_346 ? _GEN_1570 : _GEN_1538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1605 = _T_346 ? _GEN_1571 : _GEN_1539; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1606 = _T_346 ? _GEN_1572 : _GEN_1540; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1607 = _T_346 ? _GEN_1573 : _GEN_1541; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1608 = _T_346 ? _GEN_1574 : _GEN_1542; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1609 = _T_346 ? _GEN_1575 : _GEN_1543; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1610 = _T_346 ? _GEN_1576 : _GEN_1544; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1611 = _T_346 ? _GEN_1577 : _GEN_1545; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1612 = _T_346 ? _GEN_1578 : _GEN_1546; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1613 = _T_346 ? _GEN_1579 : _GEN_1547; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1614 = _T_346 ? _GEN_1580 : _GEN_1548; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1615 = _T_346 ? _GEN_1581 : _GEN_1549; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1616 = _T_346 ? _GEN_1582 : _GEN_1550; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1617 = _T_346 ? io_now_csr_mtval : _T_334; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55 194:24]
  wire  _GEN_1628 = _T_133 & _T_346; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 113:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1629 = _T_133 ? _GEN_1584 : io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1631 = _T_133 ? _GEN_1586 : _GEN_1520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1632 = _T_133 ? _GEN_1587 : _GEN_1521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1633 = _T_133 ? _GEN_1588 : _GEN_1522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1634 = _T_133 ? _GEN_1589 : _GEN_1523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1635 = _T_133 ? _GEN_1590 : _GEN_1524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1636 = _T_133 ? _GEN_1591 : _GEN_1525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1637 = _T_133 ? _GEN_1592 : _GEN_1526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1638 = _T_133 ? _GEN_1593 : _GEN_1527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1639 = _T_133 ? _GEN_1594 : _GEN_1528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1640 = _T_133 ? _GEN_1595 : _GEN_1529; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1641 = _T_133 ? _GEN_1596 : _GEN_1530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1642 = _T_133 ? _GEN_1597 : _GEN_1531; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1643 = _T_133 ? _GEN_1598 : _GEN_1532; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1644 = _T_133 ? _GEN_1599 : _GEN_1533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1645 = _T_133 ? _GEN_1600 : _GEN_1534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1646 = _T_133 ? _GEN_1601 : _GEN_1535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1647 = _T_133 ? _GEN_1602 : _GEN_1536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1648 = _T_133 ? _GEN_1603 : _GEN_1537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1649 = _T_133 ? _GEN_1604 : _GEN_1538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1650 = _T_133 ? _GEN_1605 : _GEN_1539; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1651 = _T_133 ? _GEN_1606 : _GEN_1540; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1652 = _T_133 ? _GEN_1607 : _GEN_1541; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1653 = _T_133 ? _GEN_1608 : _GEN_1542; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1654 = _T_133 ? _GEN_1609 : _GEN_1543; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1655 = _T_133 ? _GEN_1610 : _GEN_1544; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1656 = _T_133 ? _GEN_1611 : _GEN_1545; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1657 = _T_133 ? _GEN_1612 : _GEN_1546; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1658 = _T_133 ? _GEN_1613 : _GEN_1547; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1659 = _T_133 ? _GEN_1614 : _GEN_1548; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1660 = _T_133 ? _GEN_1615 : _GEN_1549; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1661 = _T_133 ? _GEN_1616 : _GEN_1550; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1662 = _T_133 ? _GEN_1617 : io_now_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1666 = 5'h1 == rd ? _next_reg_T_43 : _GEN_1631; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1667 = 5'h2 == rd ? _next_reg_T_43 : _GEN_1632; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1668 = 5'h3 == rd ? _next_reg_T_43 : _GEN_1633; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1669 = 5'h4 == rd ? _next_reg_T_43 : _GEN_1634; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1670 = 5'h5 == rd ? _next_reg_T_43 : _GEN_1635; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1671 = 5'h6 == rd ? _next_reg_T_43 : _GEN_1636; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1672 = 5'h7 == rd ? _next_reg_T_43 : _GEN_1637; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1673 = 5'h8 == rd ? _next_reg_T_43 : _GEN_1638; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1674 = 5'h9 == rd ? _next_reg_T_43 : _GEN_1639; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1675 = 5'ha == rd ? _next_reg_T_43 : _GEN_1640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1676 = 5'hb == rd ? _next_reg_T_43 : _GEN_1641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1677 = 5'hc == rd ? _next_reg_T_43 : _GEN_1642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1678 = 5'hd == rd ? _next_reg_T_43 : _GEN_1643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1679 = 5'he == rd ? _next_reg_T_43 : _GEN_1644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1680 = 5'hf == rd ? _next_reg_T_43 : _GEN_1645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1681 = 5'h10 == rd ? _next_reg_T_43 : _GEN_1646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1682 = 5'h11 == rd ? _next_reg_T_43 : _GEN_1647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1683 = 5'h12 == rd ? _next_reg_T_43 : _GEN_1648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1684 = 5'h13 == rd ? _next_reg_T_43 : _GEN_1649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1685 = 5'h14 == rd ? _next_reg_T_43 : _GEN_1650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1686 = 5'h15 == rd ? _next_reg_T_43 : _GEN_1651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1687 = 5'h16 == rd ? _next_reg_T_43 : _GEN_1652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1688 = 5'h17 == rd ? _next_reg_T_43 : _GEN_1653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1689 = 5'h18 == rd ? _next_reg_T_43 : _GEN_1654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1690 = 5'h19 == rd ? _next_reg_T_43 : _GEN_1655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1691 = 5'h1a == rd ? _next_reg_T_43 : _GEN_1656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1692 = 5'h1b == rd ? _next_reg_T_43 : _GEN_1657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1693 = 5'h1c == rd ? _next_reg_T_43 : _GEN_1658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1694 = 5'h1d == rd ? _next_reg_T_43 : _GEN_1659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1695 = 5'h1e == rd ? _next_reg_T_43 : _GEN_1660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1696 = 5'h1f == rd ? _next_reg_T_43 : _GEN_1661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire  _GEN_1697 = _T_180 | _GEN_1628; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 202:27]
  wire [63:0] _GEN_1698 = _T_180 ? _T_168 : _GEN_1629; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 203:27]
  wire [63:0] _GEN_1700 = _T_180 ? _GEN_1666 : _GEN_1631; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1701 = _T_180 ? _GEN_1667 : _GEN_1632; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1702 = _T_180 ? _GEN_1668 : _GEN_1633; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1703 = _T_180 ? _GEN_1669 : _GEN_1634; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1704 = _T_180 ? _GEN_1670 : _GEN_1635; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1705 = _T_180 ? _GEN_1671 : _GEN_1636; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1706 = _T_180 ? _GEN_1672 : _GEN_1637; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1707 = _T_180 ? _GEN_1673 : _GEN_1638; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1708 = _T_180 ? _GEN_1674 : _GEN_1639; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1709 = _T_180 ? _GEN_1675 : _GEN_1640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1710 = _T_180 ? _GEN_1676 : _GEN_1641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1711 = _T_180 ? _GEN_1677 : _GEN_1642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1712 = _T_180 ? _GEN_1678 : _GEN_1643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1713 = _T_180 ? _GEN_1679 : _GEN_1644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1714 = _T_180 ? _GEN_1680 : _GEN_1645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1715 = _T_180 ? _GEN_1681 : _GEN_1646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1716 = _T_180 ? _GEN_1682 : _GEN_1647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1717 = _T_180 ? _GEN_1683 : _GEN_1648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1718 = _T_180 ? _GEN_1684 : _GEN_1649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1719 = _T_180 ? _GEN_1685 : _GEN_1650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1720 = _T_180 ? _GEN_1686 : _GEN_1651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1721 = _T_180 ? _GEN_1687 : _GEN_1652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1722 = _T_180 ? _GEN_1688 : _GEN_1653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1723 = _T_180 ? _GEN_1689 : _GEN_1654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1724 = _T_180 ? _GEN_1690 : _GEN_1655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1725 = _T_180 ? _GEN_1691 : _GEN_1656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1726 = _T_180 ? _GEN_1692 : _GEN_1657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1727 = _T_180 ? _GEN_1693 : _GEN_1658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1728 = _T_180 ? _GEN_1694 : _GEN_1659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1729 = _T_180 ? _GEN_1695 : _GEN_1660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1730 = _T_180 ? _GEN_1696 : _GEN_1661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1731 = _T_180 ? _GEN_1662 : _T_168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 206:24]
  wire  _GEN_1741 = _T_157 ? _GEN_1697 : _GEN_1628; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1742 = _T_157 ? _GEN_1698 : _GEN_1629; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1744 = _T_157 ? _GEN_1700 : _GEN_1631; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1745 = _T_157 ? _GEN_1701 : _GEN_1632; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1746 = _T_157 ? _GEN_1702 : _GEN_1633; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1747 = _T_157 ? _GEN_1703 : _GEN_1634; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1748 = _T_157 ? _GEN_1704 : _GEN_1635; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1749 = _T_157 ? _GEN_1705 : _GEN_1636; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1750 = _T_157 ? _GEN_1706 : _GEN_1637; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1751 = _T_157 ? _GEN_1707 : _GEN_1638; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1752 = _T_157 ? _GEN_1708 : _GEN_1639; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1753 = _T_157 ? _GEN_1709 : _GEN_1640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1754 = _T_157 ? _GEN_1710 : _GEN_1641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1755 = _T_157 ? _GEN_1711 : _GEN_1642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1756 = _T_157 ? _GEN_1712 : _GEN_1643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1757 = _T_157 ? _GEN_1713 : _GEN_1644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1758 = _T_157 ? _GEN_1714 : _GEN_1645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1759 = _T_157 ? _GEN_1715 : _GEN_1646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1760 = _T_157 ? _GEN_1716 : _GEN_1647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1761 = _T_157 ? _GEN_1717 : _GEN_1648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1762 = _T_157 ? _GEN_1718 : _GEN_1649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1763 = _T_157 ? _GEN_1719 : _GEN_1650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1764 = _T_157 ? _GEN_1720 : _GEN_1651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1765 = _T_157 ? _GEN_1721 : _GEN_1652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1766 = _T_157 ? _GEN_1722 : _GEN_1653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1767 = _T_157 ? _GEN_1723 : _GEN_1654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1768 = _T_157 ? _GEN_1724 : _GEN_1655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1769 = _T_157 ? _GEN_1725 : _GEN_1656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1770 = _T_157 ? _GEN_1726 : _GEN_1657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1771 = _T_157 ? _GEN_1727 : _GEN_1658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1772 = _T_157 ? _GEN_1728 : _GEN_1659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1773 = _T_157 ? _GEN_1729 : _GEN_1660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1774 = _T_157 ? _GEN_1730 : _GEN_1661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1775 = _T_157 ? _GEN_1731 : _GEN_1662; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire  _GEN_1778 = _T_346 | _GEN_1741; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 216:29]
  wire [63:0] _GEN_1779 = _T_346 ? _T_334 : _GEN_1742; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 217:29]
  wire [63:0] _GEN_1780 = _T_346 ? _GEN_1775 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 219:26]
  wire  _GEN_1783 = _GEN_31 == _GEN_840 ? _GEN_1778 : _GEN_1741; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire [63:0] _GEN_1784 = _GEN_31 == _GEN_840 ? _GEN_1779 : _GEN_1742; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire [63:0] _GEN_1785 = _GEN_31 == _GEN_840 ? _GEN_1780 : _GEN_1775; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire  _GEN_1798 = _T_182 ? _GEN_1783 : _GEN_1741; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire [63:0] _GEN_1799 = _T_182 ? _GEN_1784 : _GEN_1742; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire [63:0] _GEN_1800 = _T_182 ? _GEN_1785 : _GEN_1775; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire  _GEN_1803 = _T_346 | _GEN_1798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 228:29]
  wire [63:0] _GEN_1804 = _T_346 ? _T_334 : _GEN_1799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 229:29]
  wire [63:0] _GEN_1805 = _T_346 ? _GEN_1800 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 231:26]
  wire  _GEN_1808 = _GEN_31 != _GEN_840 ? _GEN_1803 : _GEN_1798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire [63:0] _GEN_1809 = _GEN_31 != _GEN_840 ? _GEN_1804 : _GEN_1799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire [63:0] _GEN_1810 = _GEN_31 != _GEN_840 ? _GEN_1805 : _GEN_1800; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire  _GEN_1823 = _T_209 ? _GEN_1808 : _GEN_1798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire [63:0] _GEN_1824 = _T_209 ? _GEN_1809 : _GEN_1799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire [63:0] _GEN_1825 = _T_209 ? _GEN_1810 : _GEN_1800; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire  _GEN_1828 = _T_346 | _GEN_1823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 241:29]
  wire [63:0] _GEN_1829 = _T_346 ? _T_334 : _GEN_1824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 242:29]
  wire [63:0] _GEN_1830 = _T_346 ? _GEN_1825 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 244:26]
  wire  _GEN_1833 = $signed(_T_300) < $signed(_T_301) ? _GEN_1828 : _GEN_1823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire [63:0] _GEN_1834 = $signed(_T_300) < $signed(_T_301) ? _GEN_1829 : _GEN_1824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire [63:0] _GEN_1835 = $signed(_T_300) < $signed(_T_301) ? _GEN_1830 : _GEN_1825; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire  _GEN_1848 = _T_236 ? _GEN_1833 : _GEN_1823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire [63:0] _GEN_1849 = _T_236 ? _GEN_1834 : _GEN_1824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire [63:0] _GEN_1850 = _T_236 ? _GEN_1835 : _GEN_1825; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire  _GEN_1853 = _T_346 | _GEN_1848; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 253:29]
  wire [63:0] _GEN_1854 = _T_346 ? _T_334 : _GEN_1849; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 254:29]
  wire [63:0] _GEN_1855 = _T_346 ? _GEN_1850 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 256:26]
  wire  _GEN_1858 = _GEN_31 < _GEN_840 ? _GEN_1853 : _GEN_1848; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire [63:0] _GEN_1859 = _GEN_31 < _GEN_840 ? _GEN_1854 : _GEN_1849; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire [63:0] _GEN_1860 = _GEN_31 < _GEN_840 ? _GEN_1855 : _GEN_1850; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire  _GEN_1873 = _T_265 ? _GEN_1858 : _GEN_1848; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire [63:0] _GEN_1874 = _T_265 ? _GEN_1859 : _GEN_1849; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire [63:0] _GEN_1875 = _T_265 ? _GEN_1860 : _GEN_1850; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire  _GEN_1878 = _T_346 | _GEN_1873; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 266:29]
  wire [63:0] _GEN_1879 = _T_346 ? _T_334 : _GEN_1874; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 267:29]
  wire [63:0] _GEN_1880 = _T_346 ? _GEN_1875 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 269:26]
  wire  _GEN_1883 = $signed(_T_300) >= $signed(_T_301) ? _GEN_1878 : _GEN_1873; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire [63:0] _GEN_1884 = $signed(_T_300) >= $signed(_T_301) ? _GEN_1879 : _GEN_1874; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire [63:0] _GEN_1885 = $signed(_T_300) >= $signed(_T_301) ? _GEN_1880 : _GEN_1875; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire  _GEN_1898 = _T_292 ? _GEN_1883 : _GEN_1873; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire [63:0] _GEN_1899 = _T_292 ? _GEN_1884 : _GEN_1874; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire [63:0] _GEN_1900 = _T_292 ? _GEN_1885 : _GEN_1875; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire  _GEN_1903 = _T_346 | _GEN_1898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 278:29]
  wire [63:0] _GEN_1904 = _T_346 ? _T_334 : _GEN_1899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 279:29]
  wire [63:0] _GEN_1905 = _T_346 ? _GEN_1900 : _T_334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 281:26]
  wire  _GEN_1908 = _GEN_31 >= _GEN_840 ? _GEN_1903 : _GEN_1898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire [63:0] _GEN_1909 = _GEN_31 >= _GEN_840 ? _GEN_1904 : _GEN_1899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire [63:0] _GEN_1910 = _GEN_31 >= _GEN_840 ? _GEN_1905 : _GEN_1900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire  _GEN_1923 = _T_321 ? _GEN_1908 : _GEN_1898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire [63:0] _GEN_1924 = _T_321 ? _GEN_1909 : _GEN_1899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire [63:0] _GEN_1925 = _T_321 ? _GEN_1910 : _GEN_1900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire [5:0] next_reg_rOff = {_T_663[2:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:48]
  wire [63:0] _next_reg_T_48 = io_mem_read_data >> next_reg_rOff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:22]
  wire [63:0] _next_reg_T_49 = _next_reg_T_48 & 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire  next_reg_signBit = _next_reg_T_49[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [55:0] _next_reg_T_52 = next_reg_signBit ? 56'hffffffffffffff : 56'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_53 = {_next_reg_T_52,_next_reg_T_49[7:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_1929 = 5'h1 == rd ? _next_reg_T_53 : _GEN_1744; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1930 = 5'h2 == rd ? _next_reg_T_53 : _GEN_1745; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1931 = 5'h3 == rd ? _next_reg_T_53 : _GEN_1746; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1932 = 5'h4 == rd ? _next_reg_T_53 : _GEN_1747; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1933 = 5'h5 == rd ? _next_reg_T_53 : _GEN_1748; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1934 = 5'h6 == rd ? _next_reg_T_53 : _GEN_1749; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1935 = 5'h7 == rd ? _next_reg_T_53 : _GEN_1750; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1936 = 5'h8 == rd ? _next_reg_T_53 : _GEN_1751; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1937 = 5'h9 == rd ? _next_reg_T_53 : _GEN_1752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1938 = 5'ha == rd ? _next_reg_T_53 : _GEN_1753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1939 = 5'hb == rd ? _next_reg_T_53 : _GEN_1754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1940 = 5'hc == rd ? _next_reg_T_53 : _GEN_1755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1941 = 5'hd == rd ? _next_reg_T_53 : _GEN_1756; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1942 = 5'he == rd ? _next_reg_T_53 : _GEN_1757; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1943 = 5'hf == rd ? _next_reg_T_53 : _GEN_1758; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1944 = 5'h10 == rd ? _next_reg_T_53 : _GEN_1759; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1945 = 5'h11 == rd ? _next_reg_T_53 : _GEN_1760; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1946 = 5'h12 == rd ? _next_reg_T_53 : _GEN_1761; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1947 = 5'h13 == rd ? _next_reg_T_53 : _GEN_1762; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1948 = 5'h14 == rd ? _next_reg_T_53 : _GEN_1763; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1949 = 5'h15 == rd ? _next_reg_T_53 : _GEN_1764; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1950 = 5'h16 == rd ? _next_reg_T_53 : _GEN_1765; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1951 = 5'h17 == rd ? _next_reg_T_53 : _GEN_1766; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1952 = 5'h18 == rd ? _next_reg_T_53 : _GEN_1767; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1953 = 5'h19 == rd ? _next_reg_T_53 : _GEN_1768; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1954 = 5'h1a == rd ? _next_reg_T_53 : _GEN_1769; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1955 = 5'h1b == rd ? _next_reg_T_53 : _GEN_1770; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1956 = 5'h1c == rd ? _next_reg_T_53 : _GEN_1771; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1957 = 5'h1d == rd ? _next_reg_T_53 : _GEN_1772; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1958 = 5'h1e == rd ? _next_reg_T_53 : _GEN_1773; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_1959 = 5'h1f == rd ? _next_reg_T_53 : _GEN_1774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2005 = _T_348 ? _T_663 : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [6:0] _GEN_2006 = _T_348 ? 7'h8 : 7'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [63:0] _GEN_2008 = _T_348 ? _GEN_1929 : _GEN_1744; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2009 = _T_348 ? _GEN_1930 : _GEN_1745; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2010 = _T_348 ? _GEN_1931 : _GEN_1746; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2011 = _T_348 ? _GEN_1932 : _GEN_1747; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2012 = _T_348 ? _GEN_1933 : _GEN_1748; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2013 = _T_348 ? _GEN_1934 : _GEN_1749; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2014 = _T_348 ? _GEN_1935 : _GEN_1750; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2015 = _T_348 ? _GEN_1936 : _GEN_1751; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2016 = _T_348 ? _GEN_1937 : _GEN_1752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2017 = _T_348 ? _GEN_1938 : _GEN_1753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2018 = _T_348 ? _GEN_1939 : _GEN_1754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2019 = _T_348 ? _GEN_1940 : _GEN_1755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2020 = _T_348 ? _GEN_1941 : _GEN_1756; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2021 = _T_348 ? _GEN_1942 : _GEN_1757; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2022 = _T_348 ? _GEN_1943 : _GEN_1758; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2023 = _T_348 ? _GEN_1944 : _GEN_1759; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2024 = _T_348 ? _GEN_1945 : _GEN_1760; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2025 = _T_348 ? _GEN_1946 : _GEN_1761; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2026 = _T_348 ? _GEN_1947 : _GEN_1762; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2027 = _T_348 ? _GEN_1948 : _GEN_1763; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2028 = _T_348 ? _GEN_1949 : _GEN_1764; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2029 = _T_348 ? _GEN_1950 : _GEN_1765; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2030 = _T_348 ? _GEN_1951 : _GEN_1766; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2031 = _T_348 ? _GEN_1952 : _GEN_1767; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2032 = _T_348 ? _GEN_1953 : _GEN_1768; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2033 = _T_348 ? _GEN_1954 : _GEN_1769; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2034 = _T_348 ? _GEN_1955 : _GEN_1770; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2035 = _T_348 ? _GEN_1956 : _GEN_1771; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2036 = _T_348 ? _GEN_1957 : _GEN_1772; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2037 = _T_348 ? _GEN_1958 : _GEN_1773; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2038 = _T_348 ? _GEN_1959 : _GEN_1774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _next_reg_T_57 = _next_reg_T_48 & 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire  next_reg_signBit_1 = _next_reg_T_57[15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [47:0] _next_reg_T_60 = next_reg_signBit_1 ? 48'hffffffffffff : 48'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_61 = {_next_reg_T_60,_next_reg_T_57[15:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_2042 = 5'h1 == rd ? _next_reg_T_61 : _GEN_2008; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2043 = 5'h2 == rd ? _next_reg_T_61 : _GEN_2009; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2044 = 5'h3 == rd ? _next_reg_T_61 : _GEN_2010; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2045 = 5'h4 == rd ? _next_reg_T_61 : _GEN_2011; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2046 = 5'h5 == rd ? _next_reg_T_61 : _GEN_2012; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2047 = 5'h6 == rd ? _next_reg_T_61 : _GEN_2013; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2048 = 5'h7 == rd ? _next_reg_T_61 : _GEN_2014; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2049 = 5'h8 == rd ? _next_reg_T_61 : _GEN_2015; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2050 = 5'h9 == rd ? _next_reg_T_61 : _GEN_2016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2051 = 5'ha == rd ? _next_reg_T_61 : _GEN_2017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2052 = 5'hb == rd ? _next_reg_T_61 : _GEN_2018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2053 = 5'hc == rd ? _next_reg_T_61 : _GEN_2019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2054 = 5'hd == rd ? _next_reg_T_61 : _GEN_2020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2055 = 5'he == rd ? _next_reg_T_61 : _GEN_2021; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2056 = 5'hf == rd ? _next_reg_T_61 : _GEN_2022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2057 = 5'h10 == rd ? _next_reg_T_61 : _GEN_2023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2058 = 5'h11 == rd ? _next_reg_T_61 : _GEN_2024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2059 = 5'h12 == rd ? _next_reg_T_61 : _GEN_2025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2060 = 5'h13 == rd ? _next_reg_T_61 : _GEN_2026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2061 = 5'h14 == rd ? _next_reg_T_61 : _GEN_2027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2062 = 5'h15 == rd ? _next_reg_T_61 : _GEN_2028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2063 = 5'h16 == rd ? _next_reg_T_61 : _GEN_2029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2064 = 5'h17 == rd ? _next_reg_T_61 : _GEN_2030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2065 = 5'h18 == rd ? _next_reg_T_61 : _GEN_2031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2066 = 5'h19 == rd ? _next_reg_T_61 : _GEN_2032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2067 = 5'h1a == rd ? _next_reg_T_61 : _GEN_2033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2068 = 5'h1b == rd ? _next_reg_T_61 : _GEN_2034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2069 = 5'h1c == rd ? _next_reg_T_61 : _GEN_2035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2070 = 5'h1d == rd ? _next_reg_T_61 : _GEN_2036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2071 = 5'h1e == rd ? _next_reg_T_61 : _GEN_2037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2072 = 5'h1f == rd ? _next_reg_T_61 : _GEN_2038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire  _GEN_2073 = _T_665 | _T_348; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [63:0] _GEN_2074 = _T_665 ? _T_663 : _T_663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 303:23 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [6:0] _GEN_2075 = _T_665 ? 7'h10 : _GEN_2006; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [63:0] _GEN_2077 = _T_665 ? _GEN_2042 : _GEN_2008; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2078 = _T_665 ? _GEN_2043 : _GEN_2009; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2079 = _T_665 ? _GEN_2044 : _GEN_2010; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2080 = _T_665 ? _GEN_2045 : _GEN_2011; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2081 = _T_665 ? _GEN_2046 : _GEN_2012; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2082 = _T_665 ? _GEN_2047 : _GEN_2013; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2083 = _T_665 ? _GEN_2048 : _GEN_2014; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2084 = _T_665 ? _GEN_2049 : _GEN_2015; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2085 = _T_665 ? _GEN_2050 : _GEN_2016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2086 = _T_665 ? _GEN_2051 : _GEN_2017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2087 = _T_665 ? _GEN_2052 : _GEN_2018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2088 = _T_665 ? _GEN_2053 : _GEN_2019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2089 = _T_665 ? _GEN_2054 : _GEN_2020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2090 = _T_665 ? _GEN_2055 : _GEN_2021; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2091 = _T_665 ? _GEN_2056 : _GEN_2022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2092 = _T_665 ? _GEN_2057 : _GEN_2023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2093 = _T_665 ? _GEN_2058 : _GEN_2024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2094 = _T_665 ? _GEN_2059 : _GEN_2025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2095 = _T_665 ? _GEN_2060 : _GEN_2026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2096 = _T_665 ? _GEN_2061 : _GEN_2027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2097 = _T_665 ? _GEN_2062 : _GEN_2028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2098 = _T_665 ? _GEN_2063 : _GEN_2029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2099 = _T_665 ? _GEN_2064 : _GEN_2030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2100 = _T_665 ? _GEN_2065 : _GEN_2031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2101 = _T_665 ? _GEN_2066 : _GEN_2032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2102 = _T_665 ? _GEN_2067 : _GEN_2033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2103 = _T_665 ? _GEN_2068 : _GEN_2034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2104 = _T_665 ? _GEN_2069 : _GEN_2035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2105 = _T_665 ? _GEN_2070 : _GEN_2036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2106 = _T_665 ? _GEN_2071 : _GEN_2037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2107 = _T_665 ? _GEN_2072 : _GEN_2038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire  _GEN_2109 = _T_665 ? _GEN_1926 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_2117 = _T_368 ? _GEN_2073 : _T_348; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2118 = _T_368 ? _GEN_2074 : _GEN_2005; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [6:0] _GEN_2119 = _T_368 ? _GEN_2075 : _GEN_2006; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2121 = _T_368 ? _GEN_2077 : _GEN_2008; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2122 = _T_368 ? _GEN_2078 : _GEN_2009; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2123 = _T_368 ? _GEN_2079 : _GEN_2010; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2124 = _T_368 ? _GEN_2080 : _GEN_2011; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2125 = _T_368 ? _GEN_2081 : _GEN_2012; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2126 = _T_368 ? _GEN_2082 : _GEN_2013; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2127 = _T_368 ? _GEN_2083 : _GEN_2014; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2128 = _T_368 ? _GEN_2084 : _GEN_2015; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2129 = _T_368 ? _GEN_2085 : _GEN_2016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2130 = _T_368 ? _GEN_2086 : _GEN_2017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2131 = _T_368 ? _GEN_2087 : _GEN_2018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2132 = _T_368 ? _GEN_2088 : _GEN_2019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2133 = _T_368 ? _GEN_2089 : _GEN_2020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2134 = _T_368 ? _GEN_2090 : _GEN_2021; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2135 = _T_368 ? _GEN_2091 : _GEN_2022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2136 = _T_368 ? _GEN_2092 : _GEN_2023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2137 = _T_368 ? _GEN_2093 : _GEN_2024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2138 = _T_368 ? _GEN_2094 : _GEN_2025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2139 = _T_368 ? _GEN_2095 : _GEN_2026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2140 = _T_368 ? _GEN_2096 : _GEN_2027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2141 = _T_368 ? _GEN_2097 : _GEN_2028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2142 = _T_368 ? _GEN_2098 : _GEN_2029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2143 = _T_368 ? _GEN_2099 : _GEN_2030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2144 = _T_368 ? _GEN_2100 : _GEN_2031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2145 = _T_368 ? _GEN_2101 : _GEN_2032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2146 = _T_368 ? _GEN_2102 : _GEN_2033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2147 = _T_368 ? _GEN_2103 : _GEN_2034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2148 = _T_368 ? _GEN_2104 : _GEN_2035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2149 = _T_368 ? _GEN_2105 : _GEN_2036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2150 = _T_368 ? _GEN_2106 : _GEN_2037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2151 = _T_368 ? _GEN_2107 : _GEN_2038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire  _GEN_2153 = _T_368 ? _GEN_2109 : _GEN_1926; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _next_reg_T_65 = _next_reg_T_48 & 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire  next_reg_signBit_2 = _next_reg_T_65[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_68 = next_reg_signBit_2 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_69 = {_next_reg_T_68,_next_reg_T_65[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_2155 = 5'h1 == rd ? _next_reg_T_69 : _GEN_2121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2156 = 5'h2 == rd ? _next_reg_T_69 : _GEN_2122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2157 = 5'h3 == rd ? _next_reg_T_69 : _GEN_2123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2158 = 5'h4 == rd ? _next_reg_T_69 : _GEN_2124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2159 = 5'h5 == rd ? _next_reg_T_69 : _GEN_2125; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2160 = 5'h6 == rd ? _next_reg_T_69 : _GEN_2126; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2161 = 5'h7 == rd ? _next_reg_T_69 : _GEN_2127; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2162 = 5'h8 == rd ? _next_reg_T_69 : _GEN_2128; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2163 = 5'h9 == rd ? _next_reg_T_69 : _GEN_2129; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2164 = 5'ha == rd ? _next_reg_T_69 : _GEN_2130; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2165 = 5'hb == rd ? _next_reg_T_69 : _GEN_2131; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2166 = 5'hc == rd ? _next_reg_T_69 : _GEN_2132; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2167 = 5'hd == rd ? _next_reg_T_69 : _GEN_2133; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2168 = 5'he == rd ? _next_reg_T_69 : _GEN_2134; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2169 = 5'hf == rd ? _next_reg_T_69 : _GEN_2135; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2170 = 5'h10 == rd ? _next_reg_T_69 : _GEN_2136; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2171 = 5'h11 == rd ? _next_reg_T_69 : _GEN_2137; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2172 = 5'h12 == rd ? _next_reg_T_69 : _GEN_2138; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2173 = 5'h13 == rd ? _next_reg_T_69 : _GEN_2139; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2174 = 5'h14 == rd ? _next_reg_T_69 : _GEN_2140; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2175 = 5'h15 == rd ? _next_reg_T_69 : _GEN_2141; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2176 = 5'h16 == rd ? _next_reg_T_69 : _GEN_2142; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2177 = 5'h17 == rd ? _next_reg_T_69 : _GEN_2143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2178 = 5'h18 == rd ? _next_reg_T_69 : _GEN_2144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2179 = 5'h19 == rd ? _next_reg_T_69 : _GEN_2145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2180 = 5'h1a == rd ? _next_reg_T_69 : _GEN_2146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2181 = 5'h1b == rd ? _next_reg_T_69 : _GEN_2147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2182 = 5'h1c == rd ? _next_reg_T_69 : _GEN_2148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2183 = 5'h1d == rd ? _next_reg_T_69 : _GEN_2149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2184 = 5'h1e == rd ? _next_reg_T_69 : _GEN_2150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2185 = 5'h1f == rd ? _next_reg_T_69 : _GEN_2151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire  _GEN_2186 = _T_667 | _GEN_2117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [63:0] _GEN_2187 = _T_667 ? _T_663 : _T_663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 312:23 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [6:0] _GEN_2188 = _T_667 ? 7'h20 : _GEN_2119; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [63:0] _GEN_2190 = _T_667 ? _GEN_2155 : _GEN_2121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2191 = _T_667 ? _GEN_2156 : _GEN_2122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2192 = _T_667 ? _GEN_2157 : _GEN_2123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2193 = _T_667 ? _GEN_2158 : _GEN_2124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2194 = _T_667 ? _GEN_2159 : _GEN_2125; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2195 = _T_667 ? _GEN_2160 : _GEN_2126; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2196 = _T_667 ? _GEN_2161 : _GEN_2127; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2197 = _T_667 ? _GEN_2162 : _GEN_2128; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2198 = _T_667 ? _GEN_2163 : _GEN_2129; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2199 = _T_667 ? _GEN_2164 : _GEN_2130; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2200 = _T_667 ? _GEN_2165 : _GEN_2131; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2201 = _T_667 ? _GEN_2166 : _GEN_2132; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2202 = _T_667 ? _GEN_2167 : _GEN_2133; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2203 = _T_667 ? _GEN_2168 : _GEN_2134; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2204 = _T_667 ? _GEN_2169 : _GEN_2135; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2205 = _T_667 ? _GEN_2170 : _GEN_2136; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2206 = _T_667 ? _GEN_2171 : _GEN_2137; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2207 = _T_667 ? _GEN_2172 : _GEN_2138; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2208 = _T_667 ? _GEN_2173 : _GEN_2139; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2209 = _T_667 ? _GEN_2174 : _GEN_2140; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2210 = _T_667 ? _GEN_2175 : _GEN_2141; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2211 = _T_667 ? _GEN_2176 : _GEN_2142; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2212 = _T_667 ? _GEN_2177 : _GEN_2143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2213 = _T_667 ? _GEN_2178 : _GEN_2144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2214 = _T_667 ? _GEN_2179 : _GEN_2145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2215 = _T_667 ? _GEN_2180 : _GEN_2146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2216 = _T_667 ? _GEN_2181 : _GEN_2147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2217 = _T_667 ? _GEN_2182 : _GEN_2148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2218 = _T_667 ? _GEN_2183 : _GEN_2149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2219 = _T_667 ? _GEN_2184 : _GEN_2150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2220 = _T_667 ? _GEN_2185 : _GEN_2151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire  _GEN_2222 = _T_667 ? _GEN_2153 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_2230 = _T_388 ? _GEN_2186 : _GEN_2117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2231 = _T_388 ? _GEN_2187 : _GEN_2118; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [6:0] _GEN_2232 = _T_388 ? _GEN_2188 : _GEN_2119; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2234 = _T_388 ? _GEN_2190 : _GEN_2121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2235 = _T_388 ? _GEN_2191 : _GEN_2122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2236 = _T_388 ? _GEN_2192 : _GEN_2123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2237 = _T_388 ? _GEN_2193 : _GEN_2124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2238 = _T_388 ? _GEN_2194 : _GEN_2125; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2239 = _T_388 ? _GEN_2195 : _GEN_2126; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2240 = _T_388 ? _GEN_2196 : _GEN_2127; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2241 = _T_388 ? _GEN_2197 : _GEN_2128; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2242 = _T_388 ? _GEN_2198 : _GEN_2129; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2243 = _T_388 ? _GEN_2199 : _GEN_2130; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2244 = _T_388 ? _GEN_2200 : _GEN_2131; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2245 = _T_388 ? _GEN_2201 : _GEN_2132; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2246 = _T_388 ? _GEN_2202 : _GEN_2133; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2247 = _T_388 ? _GEN_2203 : _GEN_2134; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2248 = _T_388 ? _GEN_2204 : _GEN_2135; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2249 = _T_388 ? _GEN_2205 : _GEN_2136; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2250 = _T_388 ? _GEN_2206 : _GEN_2137; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2251 = _T_388 ? _GEN_2207 : _GEN_2138; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2252 = _T_388 ? _GEN_2208 : _GEN_2139; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2253 = _T_388 ? _GEN_2209 : _GEN_2140; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2254 = _T_388 ? _GEN_2210 : _GEN_2141; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2255 = _T_388 ? _GEN_2211 : _GEN_2142; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2256 = _T_388 ? _GEN_2212 : _GEN_2143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2257 = _T_388 ? _GEN_2213 : _GEN_2144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2258 = _T_388 ? _GEN_2214 : _GEN_2145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2259 = _T_388 ? _GEN_2215 : _GEN_2146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2260 = _T_388 ? _GEN_2216 : _GEN_2147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2261 = _T_388 ? _GEN_2217 : _GEN_2148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2262 = _T_388 ? _GEN_2218 : _GEN_2149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2263 = _T_388 ? _GEN_2219 : _GEN_2150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2264 = _T_388 ? _GEN_2220 : _GEN_2151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2266 = _T_388 ? _GEN_2222 : _GEN_2153; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _next_reg_T_75 = {56'h0,_next_reg_T_49[7:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [63:0] _GEN_2270 = 5'h1 == rd ? _next_reg_T_75 : _GEN_2234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2271 = 5'h2 == rd ? _next_reg_T_75 : _GEN_2235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2272 = 5'h3 == rd ? _next_reg_T_75 : _GEN_2236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2273 = 5'h4 == rd ? _next_reg_T_75 : _GEN_2237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2274 = 5'h5 == rd ? _next_reg_T_75 : _GEN_2238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2275 = 5'h6 == rd ? _next_reg_T_75 : _GEN_2239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2276 = 5'h7 == rd ? _next_reg_T_75 : _GEN_2240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2277 = 5'h8 == rd ? _next_reg_T_75 : _GEN_2241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2278 = 5'h9 == rd ? _next_reg_T_75 : _GEN_2242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2279 = 5'ha == rd ? _next_reg_T_75 : _GEN_2243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2280 = 5'hb == rd ? _next_reg_T_75 : _GEN_2244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2281 = 5'hc == rd ? _next_reg_T_75 : _GEN_2245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2282 = 5'hd == rd ? _next_reg_T_75 : _GEN_2246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2283 = 5'he == rd ? _next_reg_T_75 : _GEN_2247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2284 = 5'hf == rd ? _next_reg_T_75 : _GEN_2248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2285 = 5'h10 == rd ? _next_reg_T_75 : _GEN_2249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2286 = 5'h11 == rd ? _next_reg_T_75 : _GEN_2250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2287 = 5'h12 == rd ? _next_reg_T_75 : _GEN_2251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2288 = 5'h13 == rd ? _next_reg_T_75 : _GEN_2252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2289 = 5'h14 == rd ? _next_reg_T_75 : _GEN_2253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2290 = 5'h15 == rd ? _next_reg_T_75 : _GEN_2254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2291 = 5'h16 == rd ? _next_reg_T_75 : _GEN_2255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2292 = 5'h17 == rd ? _next_reg_T_75 : _GEN_2256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2293 = 5'h18 == rd ? _next_reg_T_75 : _GEN_2257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2294 = 5'h19 == rd ? _next_reg_T_75 : _GEN_2258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2295 = 5'h1a == rd ? _next_reg_T_75 : _GEN_2259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2296 = 5'h1b == rd ? _next_reg_T_75 : _GEN_2260; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2297 = 5'h1c == rd ? _next_reg_T_75 : _GEN_2261; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2298 = 5'h1d == rd ? _next_reg_T_75 : _GEN_2262; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2299 = 5'h1e == rd ? _next_reg_T_75 : _GEN_2263; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2300 = 5'h1f == rd ? _next_reg_T_75 : _GEN_2264; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire  _GEN_2310 = _T_408 | _GEN_2230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [63:0] _GEN_2311 = _T_408 ? _T_663 : _GEN_2231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [6:0] _GEN_2312 = _T_408 ? 7'h8 : _GEN_2232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [63:0] _GEN_2314 = _T_408 ? _GEN_2270 : _GEN_2234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2315 = _T_408 ? _GEN_2271 : _GEN_2235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2316 = _T_408 ? _GEN_2272 : _GEN_2236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2317 = _T_408 ? _GEN_2273 : _GEN_2237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2318 = _T_408 ? _GEN_2274 : _GEN_2238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2319 = _T_408 ? _GEN_2275 : _GEN_2239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2320 = _T_408 ? _GEN_2276 : _GEN_2240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2321 = _T_408 ? _GEN_2277 : _GEN_2241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2322 = _T_408 ? _GEN_2278 : _GEN_2242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2323 = _T_408 ? _GEN_2279 : _GEN_2243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2324 = _T_408 ? _GEN_2280 : _GEN_2244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2325 = _T_408 ? _GEN_2281 : _GEN_2245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2326 = _T_408 ? _GEN_2282 : _GEN_2246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2327 = _T_408 ? _GEN_2283 : _GEN_2247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2328 = _T_408 ? _GEN_2284 : _GEN_2248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2329 = _T_408 ? _GEN_2285 : _GEN_2249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2330 = _T_408 ? _GEN_2286 : _GEN_2250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2331 = _T_408 ? _GEN_2287 : _GEN_2251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2332 = _T_408 ? _GEN_2288 : _GEN_2252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2333 = _T_408 ? _GEN_2289 : _GEN_2253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2334 = _T_408 ? _GEN_2290 : _GEN_2254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2335 = _T_408 ? _GEN_2291 : _GEN_2255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2336 = _T_408 ? _GEN_2292 : _GEN_2256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2337 = _T_408 ? _GEN_2293 : _GEN_2257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2338 = _T_408 ? _GEN_2294 : _GEN_2258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2339 = _T_408 ? _GEN_2295 : _GEN_2259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2340 = _T_408 ? _GEN_2296 : _GEN_2260; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2341 = _T_408 ? _GEN_2297 : _GEN_2261; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2342 = _T_408 ? _GEN_2298 : _GEN_2262; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2343 = _T_408 ? _GEN_2299 : _GEN_2263; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2344 = _T_408 ? _GEN_2300 : _GEN_2264; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _next_reg_T_81 = {48'h0,_next_reg_T_57[15:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [63:0] _GEN_2346 = 5'h1 == rd ? _next_reg_T_81 : _GEN_2314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2347 = 5'h2 == rd ? _next_reg_T_81 : _GEN_2315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2348 = 5'h3 == rd ? _next_reg_T_81 : _GEN_2316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2349 = 5'h4 == rd ? _next_reg_T_81 : _GEN_2317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2350 = 5'h5 == rd ? _next_reg_T_81 : _GEN_2318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2351 = 5'h6 == rd ? _next_reg_T_81 : _GEN_2319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2352 = 5'h7 == rd ? _next_reg_T_81 : _GEN_2320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2353 = 5'h8 == rd ? _next_reg_T_81 : _GEN_2321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2354 = 5'h9 == rd ? _next_reg_T_81 : _GEN_2322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2355 = 5'ha == rd ? _next_reg_T_81 : _GEN_2323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2356 = 5'hb == rd ? _next_reg_T_81 : _GEN_2324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2357 = 5'hc == rd ? _next_reg_T_81 : _GEN_2325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2358 = 5'hd == rd ? _next_reg_T_81 : _GEN_2326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2359 = 5'he == rd ? _next_reg_T_81 : _GEN_2327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2360 = 5'hf == rd ? _next_reg_T_81 : _GEN_2328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2361 = 5'h10 == rd ? _next_reg_T_81 : _GEN_2329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2362 = 5'h11 == rd ? _next_reg_T_81 : _GEN_2330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2363 = 5'h12 == rd ? _next_reg_T_81 : _GEN_2331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2364 = 5'h13 == rd ? _next_reg_T_81 : _GEN_2332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2365 = 5'h14 == rd ? _next_reg_T_81 : _GEN_2333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2366 = 5'h15 == rd ? _next_reg_T_81 : _GEN_2334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2367 = 5'h16 == rd ? _next_reg_T_81 : _GEN_2335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2368 = 5'h17 == rd ? _next_reg_T_81 : _GEN_2336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2369 = 5'h18 == rd ? _next_reg_T_81 : _GEN_2337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2370 = 5'h19 == rd ? _next_reg_T_81 : _GEN_2338; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2371 = 5'h1a == rd ? _next_reg_T_81 : _GEN_2339; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2372 = 5'h1b == rd ? _next_reg_T_81 : _GEN_2340; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2373 = 5'h1c == rd ? _next_reg_T_81 : _GEN_2341; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2374 = 5'h1d == rd ? _next_reg_T_81 : _GEN_2342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2375 = 5'h1e == rd ? _next_reg_T_81 : _GEN_2343; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_2376 = 5'h1f == rd ? _next_reg_T_81 : _GEN_2344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire  _GEN_2377 = _T_665 | _GEN_2310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [6:0] _GEN_2379 = _T_665 ? 7'h10 : _GEN_2312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [63:0] _GEN_2381 = _T_665 ? _GEN_2346 : _GEN_2314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2382 = _T_665 ? _GEN_2347 : _GEN_2315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2383 = _T_665 ? _GEN_2348 : _GEN_2316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2384 = _T_665 ? _GEN_2349 : _GEN_2317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2385 = _T_665 ? _GEN_2350 : _GEN_2318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2386 = _T_665 ? _GEN_2351 : _GEN_2319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2387 = _T_665 ? _GEN_2352 : _GEN_2320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2388 = _T_665 ? _GEN_2353 : _GEN_2321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2389 = _T_665 ? _GEN_2354 : _GEN_2322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2390 = _T_665 ? _GEN_2355 : _GEN_2323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2391 = _T_665 ? _GEN_2356 : _GEN_2324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2392 = _T_665 ? _GEN_2357 : _GEN_2325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2393 = _T_665 ? _GEN_2358 : _GEN_2326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2394 = _T_665 ? _GEN_2359 : _GEN_2327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2395 = _T_665 ? _GEN_2360 : _GEN_2328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2396 = _T_665 ? _GEN_2361 : _GEN_2329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2397 = _T_665 ? _GEN_2362 : _GEN_2330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2398 = _T_665 ? _GEN_2363 : _GEN_2331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2399 = _T_665 ? _GEN_2364 : _GEN_2332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2400 = _T_665 ? _GEN_2365 : _GEN_2333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2401 = _T_665 ? _GEN_2366 : _GEN_2334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2402 = _T_665 ? _GEN_2367 : _GEN_2335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2403 = _T_665 ? _GEN_2368 : _GEN_2336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2404 = _T_665 ? _GEN_2369 : _GEN_2337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2405 = _T_665 ? _GEN_2370 : _GEN_2338; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2406 = _T_665 ? _GEN_2371 : _GEN_2339; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2407 = _T_665 ? _GEN_2372 : _GEN_2340; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2408 = _T_665 ? _GEN_2373 : _GEN_2341; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2409 = _T_665 ? _GEN_2374 : _GEN_2342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2410 = _T_665 ? _GEN_2375 : _GEN_2343; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_2411 = _T_665 ? _GEN_2376 : _GEN_2344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire  _GEN_2413 = _T_665 ? _GEN_2266 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_2421 = _T_427 ? _GEN_2377 : _GEN_2310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2422 = _T_427 ? _GEN_2074 : _GEN_2311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [6:0] _GEN_2423 = _T_427 ? _GEN_2379 : _GEN_2312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2425 = _T_427 ? _GEN_2381 : _GEN_2314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2426 = _T_427 ? _GEN_2382 : _GEN_2315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2427 = _T_427 ? _GEN_2383 : _GEN_2316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2428 = _T_427 ? _GEN_2384 : _GEN_2317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2429 = _T_427 ? _GEN_2385 : _GEN_2318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2430 = _T_427 ? _GEN_2386 : _GEN_2319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2431 = _T_427 ? _GEN_2387 : _GEN_2320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2432 = _T_427 ? _GEN_2388 : _GEN_2321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2433 = _T_427 ? _GEN_2389 : _GEN_2322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2434 = _T_427 ? _GEN_2390 : _GEN_2323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2435 = _T_427 ? _GEN_2391 : _GEN_2324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2436 = _T_427 ? _GEN_2392 : _GEN_2325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2437 = _T_427 ? _GEN_2393 : _GEN_2326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2438 = _T_427 ? _GEN_2394 : _GEN_2327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2439 = _T_427 ? _GEN_2395 : _GEN_2328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2440 = _T_427 ? _GEN_2396 : _GEN_2329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2441 = _T_427 ? _GEN_2397 : _GEN_2330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2442 = _T_427 ? _GEN_2398 : _GEN_2331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2443 = _T_427 ? _GEN_2399 : _GEN_2332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2444 = _T_427 ? _GEN_2400 : _GEN_2333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2445 = _T_427 ? _GEN_2401 : _GEN_2334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2446 = _T_427 ? _GEN_2402 : _GEN_2335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2447 = _T_427 ? _GEN_2403 : _GEN_2336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2448 = _T_427 ? _GEN_2404 : _GEN_2337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2449 = _T_427 ? _GEN_2405 : _GEN_2338; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2450 = _T_427 ? _GEN_2406 : _GEN_2339; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2451 = _T_427 ? _GEN_2407 : _GEN_2340; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2452 = _T_427 ? _GEN_2408 : _GEN_2341; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2453 = _T_427 ? _GEN_2409 : _GEN_2342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2454 = _T_427 ? _GEN_2410 : _GEN_2343; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2455 = _T_427 ? _GEN_2411 : _GEN_2344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire  _GEN_2457 = _T_427 ? _GEN_2413 : _GEN_2266; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_2471 = _T_447 ? _T_663 : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/LoadStore.scala 83:26 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [6:0] _GEN_2472 = _T_447 ? 7'h8 : 7'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/LoadStore.scala 84:26 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [63:0] _GEN_2473 = _T_447 ? {{56'd0}, _GEN_840[7:0]} : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:26 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire  _GEN_2474 = _T_665 | _T_447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 82:26]
  wire [6:0] _GEN_2476 = _T_665 ? 7'h10 : _GEN_2472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 84:26]
  wire [63:0] _GEN_2477 = _T_665 ? {{48'd0}, _GEN_840[15:0]} : _GEN_2473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:26]
  wire  _GEN_2479 = _T_665 ? _GEN_2457 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_2488 = _T_470 ? _GEN_2474 : _T_447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [63:0] _GEN_2489 = _T_470 ? _GEN_2074 : _GEN_2471; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [6:0] _GEN_2490 = _T_470 ? _GEN_2476 : _GEN_2472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [63:0] _GEN_2491 = _T_470 ? _GEN_2477 : _GEN_2473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire  _GEN_2493 = _T_470 ? _GEN_2479 : _GEN_2457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire  _GEN_2494 = _T_667 | _GEN_2488; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 82:26]
  wire [6:0] _GEN_2496 = _T_667 ? 7'h20 : _GEN_2490; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 84:26]
  wire [63:0] _GEN_2497 = _T_667 ? {{32'd0}, _GEN_840[31:0]} : _GEN_2491; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:26]
  wire  _GEN_2499 = _T_667 ? _GEN_2493 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_2508 = _T_494 ? _GEN_2494 : _GEN_2488; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [63:0] _GEN_2509 = _T_494 ? _GEN_2187 : _GEN_2489; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [6:0] _GEN_2510 = _T_494 ? _GEN_2496 : _GEN_2490; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [63:0] _GEN_2511 = _T_494 ? _GEN_2497 : _GEN_2491; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire  _GEN_2513 = _T_494 ? _GEN_2499 : _GEN_2493; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire  _GEN_2522 = _T_518 | _GEN_2513; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_2529 = 2'h3 == io_now_internal_privilegeMode | (2'h1 == io_now_internal_privilegeMode | (2'h0 ==
    io_now_internal_privilegeMode | _GEN_2522)); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_2540 = _T_524 ? _GEN_2529 : _GEN_2522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23]
  wire  next_reg_signBit_3 = _T_663[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_86 = next_reg_signBit_3 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_87 = {_next_reg_T_86,_T_663[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_2551 = 5'h1 == rd ? _next_reg_T_87 : _GEN_2425; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2552 = 5'h2 == rd ? _next_reg_T_87 : _GEN_2426; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2553 = 5'h3 == rd ? _next_reg_T_87 : _GEN_2427; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2554 = 5'h4 == rd ? _next_reg_T_87 : _GEN_2428; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2555 = 5'h5 == rd ? _next_reg_T_87 : _GEN_2429; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2556 = 5'h6 == rd ? _next_reg_T_87 : _GEN_2430; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2557 = 5'h7 == rd ? _next_reg_T_87 : _GEN_2431; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2558 = 5'h8 == rd ? _next_reg_T_87 : _GEN_2432; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2559 = 5'h9 == rd ? _next_reg_T_87 : _GEN_2433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2560 = 5'ha == rd ? _next_reg_T_87 : _GEN_2434; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2561 = 5'hb == rd ? _next_reg_T_87 : _GEN_2435; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2562 = 5'hc == rd ? _next_reg_T_87 : _GEN_2436; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2563 = 5'hd == rd ? _next_reg_T_87 : _GEN_2437; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2564 = 5'he == rd ? _next_reg_T_87 : _GEN_2438; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2565 = 5'hf == rd ? _next_reg_T_87 : _GEN_2439; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2566 = 5'h10 == rd ? _next_reg_T_87 : _GEN_2440; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2567 = 5'h11 == rd ? _next_reg_T_87 : _GEN_2441; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2568 = 5'h12 == rd ? _next_reg_T_87 : _GEN_2442; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2569 = 5'h13 == rd ? _next_reg_T_87 : _GEN_2443; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2570 = 5'h14 == rd ? _next_reg_T_87 : _GEN_2444; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2571 = 5'h15 == rd ? _next_reg_T_87 : _GEN_2445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2572 = 5'h16 == rd ? _next_reg_T_87 : _GEN_2446; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2573 = 5'h17 == rd ? _next_reg_T_87 : _GEN_2447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2574 = 5'h18 == rd ? _next_reg_T_87 : _GEN_2448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2575 = 5'h19 == rd ? _next_reg_T_87 : _GEN_2449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2576 = 5'h1a == rd ? _next_reg_T_87 : _GEN_2450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2577 = 5'h1b == rd ? _next_reg_T_87 : _GEN_2451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2578 = 5'h1c == rd ? _next_reg_T_87 : _GEN_2452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2579 = 5'h1d == rd ? _next_reg_T_87 : _GEN_2453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2580 = 5'h1e == rd ? _next_reg_T_87 : _GEN_2454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2581 = 5'h1f == rd ? _next_reg_T_87 : _GEN_2455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_2590 = _T_539 ? _GEN_2551 : _GEN_2425; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2591 = _T_539 ? _GEN_2552 : _GEN_2426; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2592 = _T_539 ? _GEN_2553 : _GEN_2427; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2593 = _T_539 ? _GEN_2554 : _GEN_2428; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2594 = _T_539 ? _GEN_2555 : _GEN_2429; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2595 = _T_539 ? _GEN_2556 : _GEN_2430; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2596 = _T_539 ? _GEN_2557 : _GEN_2431; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2597 = _T_539 ? _GEN_2558 : _GEN_2432; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2598 = _T_539 ? _GEN_2559 : _GEN_2433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2599 = _T_539 ? _GEN_2560 : _GEN_2434; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2600 = _T_539 ? _GEN_2561 : _GEN_2435; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2601 = _T_539 ? _GEN_2562 : _GEN_2436; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2602 = _T_539 ? _GEN_2563 : _GEN_2437; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2603 = _T_539 ? _GEN_2564 : _GEN_2438; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2604 = _T_539 ? _GEN_2565 : _GEN_2439; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2605 = _T_539 ? _GEN_2566 : _GEN_2440; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2606 = _T_539 ? _GEN_2567 : _GEN_2441; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2607 = _T_539 ? _GEN_2568 : _GEN_2442; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2608 = _T_539 ? _GEN_2569 : _GEN_2443; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2609 = _T_539 ? _GEN_2570 : _GEN_2444; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2610 = _T_539 ? _GEN_2571 : _GEN_2445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2611 = _T_539 ? _GEN_2572 : _GEN_2446; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2612 = _T_539 ? _GEN_2573 : _GEN_2447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2613 = _T_539 ? _GEN_2574 : _GEN_2448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2614 = _T_539 ? _GEN_2575 : _GEN_2449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2615 = _T_539 ? _GEN_2576 : _GEN_2450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2616 = _T_539 ? _GEN_2577 : _GEN_2451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2617 = _T_539 ? _GEN_2578 : _GEN_2452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2618 = _T_539 ? _GEN_2579 : _GEN_2453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2619 = _T_539 ? _GEN_2580 : _GEN_2454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_2620 = _T_539 ? _GEN_2581 : _GEN_2455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [126:0] _GEN_67 = {{63'd0}, _GEN_31}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:62]
  wire [126:0] _next_reg_T_89 = _GEN_67 << imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:62]
  wire [63:0] _GEN_2622 = 5'h1 == rd ? _next_reg_T_89[63:0] : _GEN_2590; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2623 = 5'h2 == rd ? _next_reg_T_89[63:0] : _GEN_2591; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2624 = 5'h3 == rd ? _next_reg_T_89[63:0] : _GEN_2592; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2625 = 5'h4 == rd ? _next_reg_T_89[63:0] : _GEN_2593; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2626 = 5'h5 == rd ? _next_reg_T_89[63:0] : _GEN_2594; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2627 = 5'h6 == rd ? _next_reg_T_89[63:0] : _GEN_2595; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2628 = 5'h7 == rd ? _next_reg_T_89[63:0] : _GEN_2596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2629 = 5'h8 == rd ? _next_reg_T_89[63:0] : _GEN_2597; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2630 = 5'h9 == rd ? _next_reg_T_89[63:0] : _GEN_2598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2631 = 5'ha == rd ? _next_reg_T_89[63:0] : _GEN_2599; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2632 = 5'hb == rd ? _next_reg_T_89[63:0] : _GEN_2600; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2633 = 5'hc == rd ? _next_reg_T_89[63:0] : _GEN_2601; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2634 = 5'hd == rd ? _next_reg_T_89[63:0] : _GEN_2602; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2635 = 5'he == rd ? _next_reg_T_89[63:0] : _GEN_2603; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2636 = 5'hf == rd ? _next_reg_T_89[63:0] : _GEN_2604; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2637 = 5'h10 == rd ? _next_reg_T_89[63:0] : _GEN_2605; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2638 = 5'h11 == rd ? _next_reg_T_89[63:0] : _GEN_2606; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2639 = 5'h12 == rd ? _next_reg_T_89[63:0] : _GEN_2607; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2640 = 5'h13 == rd ? _next_reg_T_89[63:0] : _GEN_2608; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2641 = 5'h14 == rd ? _next_reg_T_89[63:0] : _GEN_2609; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2642 = 5'h15 == rd ? _next_reg_T_89[63:0] : _GEN_2610; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2643 = 5'h16 == rd ? _next_reg_T_89[63:0] : _GEN_2611; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2644 = 5'h17 == rd ? _next_reg_T_89[63:0] : _GEN_2612; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2645 = 5'h18 == rd ? _next_reg_T_89[63:0] : _GEN_2613; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2646 = 5'h19 == rd ? _next_reg_T_89[63:0] : _GEN_2614; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2647 = 5'h1a == rd ? _next_reg_T_89[63:0] : _GEN_2615; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2648 = 5'h1b == rd ? _next_reg_T_89[63:0] : _GEN_2616; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2649 = 5'h1c == rd ? _next_reg_T_89[63:0] : _GEN_2617; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2650 = 5'h1d == rd ? _next_reg_T_89[63:0] : _GEN_2618; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2651 = 5'h1e == rd ? _next_reg_T_89[63:0] : _GEN_2619; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2652 = 5'h1f == rd ? _next_reg_T_89[63:0] : _GEN_2620; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_2661 = _T_545 ? _GEN_2622 : _GEN_2590; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2662 = _T_545 ? _GEN_2623 : _GEN_2591; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2663 = _T_545 ? _GEN_2624 : _GEN_2592; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2664 = _T_545 ? _GEN_2625 : _GEN_2593; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2665 = _T_545 ? _GEN_2626 : _GEN_2594; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2666 = _T_545 ? _GEN_2627 : _GEN_2595; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2667 = _T_545 ? _GEN_2628 : _GEN_2596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2668 = _T_545 ? _GEN_2629 : _GEN_2597; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2669 = _T_545 ? _GEN_2630 : _GEN_2598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2670 = _T_545 ? _GEN_2631 : _GEN_2599; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2671 = _T_545 ? _GEN_2632 : _GEN_2600; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2672 = _T_545 ? _GEN_2633 : _GEN_2601; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2673 = _T_545 ? _GEN_2634 : _GEN_2602; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2674 = _T_545 ? _GEN_2635 : _GEN_2603; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2675 = _T_545 ? _GEN_2636 : _GEN_2604; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2676 = _T_545 ? _GEN_2637 : _GEN_2605; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2677 = _T_545 ? _GEN_2638 : _GEN_2606; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2678 = _T_545 ? _GEN_2639 : _GEN_2607; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2679 = _T_545 ? _GEN_2640 : _GEN_2608; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2680 = _T_545 ? _GEN_2641 : _GEN_2609; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2681 = _T_545 ? _GEN_2642 : _GEN_2610; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2682 = _T_545 ? _GEN_2643 : _GEN_2611; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2683 = _T_545 ? _GEN_2644 : _GEN_2612; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2684 = _T_545 ? _GEN_2645 : _GEN_2613; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2685 = _T_545 ? _GEN_2646 : _GEN_2614; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2686 = _T_545 ? _GEN_2647 : _GEN_2615; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2687 = _T_545 ? _GEN_2648 : _GEN_2616; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2688 = _T_545 ? _GEN_2649 : _GEN_2617; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2689 = _T_545 ? _GEN_2650 : _GEN_2618; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2690 = _T_545 ? _GEN_2651 : _GEN_2619; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_2691 = _T_545 ? _GEN_2652 : _GEN_2620; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _next_reg_T_91 = _GEN_31 >> imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:62]
  wire [63:0] _GEN_2693 = 5'h1 == rd ? _next_reg_T_91 : _GEN_2661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2694 = 5'h2 == rd ? _next_reg_T_91 : _GEN_2662; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2695 = 5'h3 == rd ? _next_reg_T_91 : _GEN_2663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2696 = 5'h4 == rd ? _next_reg_T_91 : _GEN_2664; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2697 = 5'h5 == rd ? _next_reg_T_91 : _GEN_2665; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2698 = 5'h6 == rd ? _next_reg_T_91 : _GEN_2666; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2699 = 5'h7 == rd ? _next_reg_T_91 : _GEN_2667; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2700 = 5'h8 == rd ? _next_reg_T_91 : _GEN_2668; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2701 = 5'h9 == rd ? _next_reg_T_91 : _GEN_2669; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2702 = 5'ha == rd ? _next_reg_T_91 : _GEN_2670; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2703 = 5'hb == rd ? _next_reg_T_91 : _GEN_2671; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2704 = 5'hc == rd ? _next_reg_T_91 : _GEN_2672; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2705 = 5'hd == rd ? _next_reg_T_91 : _GEN_2673; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2706 = 5'he == rd ? _next_reg_T_91 : _GEN_2674; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2707 = 5'hf == rd ? _next_reg_T_91 : _GEN_2675; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2708 = 5'h10 == rd ? _next_reg_T_91 : _GEN_2676; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2709 = 5'h11 == rd ? _next_reg_T_91 : _GEN_2677; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2710 = 5'h12 == rd ? _next_reg_T_91 : _GEN_2678; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2711 = 5'h13 == rd ? _next_reg_T_91 : _GEN_2679; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2712 = 5'h14 == rd ? _next_reg_T_91 : _GEN_2680; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2713 = 5'h15 == rd ? _next_reg_T_91 : _GEN_2681; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2714 = 5'h16 == rd ? _next_reg_T_91 : _GEN_2682; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2715 = 5'h17 == rd ? _next_reg_T_91 : _GEN_2683; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2716 = 5'h18 == rd ? _next_reg_T_91 : _GEN_2684; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2717 = 5'h19 == rd ? _next_reg_T_91 : _GEN_2685; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2718 = 5'h1a == rd ? _next_reg_T_91 : _GEN_2686; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2719 = 5'h1b == rd ? _next_reg_T_91 : _GEN_2687; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2720 = 5'h1c == rd ? _next_reg_T_91 : _GEN_2688; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2721 = 5'h1d == rd ? _next_reg_T_91 : _GEN_2689; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2722 = 5'h1e == rd ? _next_reg_T_91 : _GEN_2690; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2723 = 5'h1f == rd ? _next_reg_T_91 : _GEN_2691; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_2732 = _T_551 ? _GEN_2693 : _GEN_2661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2733 = _T_551 ? _GEN_2694 : _GEN_2662; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2734 = _T_551 ? _GEN_2695 : _GEN_2663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2735 = _T_551 ? _GEN_2696 : _GEN_2664; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2736 = _T_551 ? _GEN_2697 : _GEN_2665; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2737 = _T_551 ? _GEN_2698 : _GEN_2666; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2738 = _T_551 ? _GEN_2699 : _GEN_2667; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2739 = _T_551 ? _GEN_2700 : _GEN_2668; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2740 = _T_551 ? _GEN_2701 : _GEN_2669; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2741 = _T_551 ? _GEN_2702 : _GEN_2670; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2742 = _T_551 ? _GEN_2703 : _GEN_2671; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2743 = _T_551 ? _GEN_2704 : _GEN_2672; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2744 = _T_551 ? _GEN_2705 : _GEN_2673; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2745 = _T_551 ? _GEN_2706 : _GEN_2674; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2746 = _T_551 ? _GEN_2707 : _GEN_2675; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2747 = _T_551 ? _GEN_2708 : _GEN_2676; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2748 = _T_551 ? _GEN_2709 : _GEN_2677; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2749 = _T_551 ? _GEN_2710 : _GEN_2678; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2750 = _T_551 ? _GEN_2711 : _GEN_2679; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2751 = _T_551 ? _GEN_2712 : _GEN_2680; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2752 = _T_551 ? _GEN_2713 : _GEN_2681; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2753 = _T_551 ? _GEN_2714 : _GEN_2682; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2754 = _T_551 ? _GEN_2715 : _GEN_2683; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2755 = _T_551 ? _GEN_2716 : _GEN_2684; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2756 = _T_551 ? _GEN_2717 : _GEN_2685; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2757 = _T_551 ? _GEN_2718 : _GEN_2686; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2758 = _T_551 ? _GEN_2719 : _GEN_2687; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2759 = _T_551 ? _GEN_2720 : _GEN_2688; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2760 = _T_551 ? _GEN_2721 : _GEN_2689; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2761 = _T_551 ? _GEN_2722 : _GEN_2690; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_2762 = _T_551 ? _GEN_2723 : _GEN_2691; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _next_reg_T_95 = $signed(_T_300) >>> imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:84]
  wire [63:0] _GEN_2764 = 5'h1 == rd ? _next_reg_T_95 : _GEN_2732; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2765 = 5'h2 == rd ? _next_reg_T_95 : _GEN_2733; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2766 = 5'h3 == rd ? _next_reg_T_95 : _GEN_2734; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2767 = 5'h4 == rd ? _next_reg_T_95 : _GEN_2735; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2768 = 5'h5 == rd ? _next_reg_T_95 : _GEN_2736; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2769 = 5'h6 == rd ? _next_reg_T_95 : _GEN_2737; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2770 = 5'h7 == rd ? _next_reg_T_95 : _GEN_2738; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2771 = 5'h8 == rd ? _next_reg_T_95 : _GEN_2739; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2772 = 5'h9 == rd ? _next_reg_T_95 : _GEN_2740; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2773 = 5'ha == rd ? _next_reg_T_95 : _GEN_2741; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2774 = 5'hb == rd ? _next_reg_T_95 : _GEN_2742; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2775 = 5'hc == rd ? _next_reg_T_95 : _GEN_2743; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2776 = 5'hd == rd ? _next_reg_T_95 : _GEN_2744; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2777 = 5'he == rd ? _next_reg_T_95 : _GEN_2745; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2778 = 5'hf == rd ? _next_reg_T_95 : _GEN_2746; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2779 = 5'h10 == rd ? _next_reg_T_95 : _GEN_2747; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2780 = 5'h11 == rd ? _next_reg_T_95 : _GEN_2748; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2781 = 5'h12 == rd ? _next_reg_T_95 : _GEN_2749; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2782 = 5'h13 == rd ? _next_reg_T_95 : _GEN_2750; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2783 = 5'h14 == rd ? _next_reg_T_95 : _GEN_2751; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2784 = 5'h15 == rd ? _next_reg_T_95 : _GEN_2752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2785 = 5'h16 == rd ? _next_reg_T_95 : _GEN_2753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2786 = 5'h17 == rd ? _next_reg_T_95 : _GEN_2754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2787 = 5'h18 == rd ? _next_reg_T_95 : _GEN_2755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2788 = 5'h19 == rd ? _next_reg_T_95 : _GEN_2756; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2789 = 5'h1a == rd ? _next_reg_T_95 : _GEN_2757; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2790 = 5'h1b == rd ? _next_reg_T_95 : _GEN_2758; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2791 = 5'h1c == rd ? _next_reg_T_95 : _GEN_2759; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2792 = 5'h1d == rd ? _next_reg_T_95 : _GEN_2760; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2793 = 5'h1e == rd ? _next_reg_T_95 : _GEN_2761; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2794 = 5'h1f == rd ? _next_reg_T_95 : _GEN_2762; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_2803 = _T_557 ? _GEN_2764 : _GEN_2732; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2804 = _T_557 ? _GEN_2765 : _GEN_2733; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2805 = _T_557 ? _GEN_2766 : _GEN_2734; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2806 = _T_557 ? _GEN_2767 : _GEN_2735; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2807 = _T_557 ? _GEN_2768 : _GEN_2736; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2808 = _T_557 ? _GEN_2769 : _GEN_2737; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2809 = _T_557 ? _GEN_2770 : _GEN_2738; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2810 = _T_557 ? _GEN_2771 : _GEN_2739; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2811 = _T_557 ? _GEN_2772 : _GEN_2740; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2812 = _T_557 ? _GEN_2773 : _GEN_2741; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2813 = _T_557 ? _GEN_2774 : _GEN_2742; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2814 = _T_557 ? _GEN_2775 : _GEN_2743; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2815 = _T_557 ? _GEN_2776 : _GEN_2744; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2816 = _T_557 ? _GEN_2777 : _GEN_2745; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2817 = _T_557 ? _GEN_2778 : _GEN_2746; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2818 = _T_557 ? _GEN_2779 : _GEN_2747; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2819 = _T_557 ? _GEN_2780 : _GEN_2748; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2820 = _T_557 ? _GEN_2781 : _GEN_2749; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2821 = _T_557 ? _GEN_2782 : _GEN_2750; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2822 = _T_557 ? _GEN_2783 : _GEN_2751; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2823 = _T_557 ? _GEN_2784 : _GEN_2752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2824 = _T_557 ? _GEN_2785 : _GEN_2753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2825 = _T_557 ? _GEN_2786 : _GEN_2754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2826 = _T_557 ? _GEN_2787 : _GEN_2755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2827 = _T_557 ? _GEN_2788 : _GEN_2756; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2828 = _T_557 ? _GEN_2789 : _GEN_2757; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2829 = _T_557 ? _GEN_2790 : _GEN_2758; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2830 = _T_557 ? _GEN_2791 : _GEN_2759; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2831 = _T_557 ? _GEN_2792 : _GEN_2760; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2832 = _T_557 ? _GEN_2793 : _GEN_2761; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_2833 = _T_557 ? _GEN_2794 : _GEN_2762; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [62:0] _GEN_69 = {{31'd0}, _GEN_31[31:0]}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:79]
  wire [62:0] _next_reg_T_98 = _GEN_69 << imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:79]
  wire  next_reg_signBit_4 = _next_reg_T_98[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_101 = next_reg_signBit_4 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_102 = {_next_reg_T_101,_next_reg_T_98[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_2835 = 5'h1 == rd ? _next_reg_T_102 : _GEN_2803; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2836 = 5'h2 == rd ? _next_reg_T_102 : _GEN_2804; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2837 = 5'h3 == rd ? _next_reg_T_102 : _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2838 = 5'h4 == rd ? _next_reg_T_102 : _GEN_2806; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2839 = 5'h5 == rd ? _next_reg_T_102 : _GEN_2807; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2840 = 5'h6 == rd ? _next_reg_T_102 : _GEN_2808; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2841 = 5'h7 == rd ? _next_reg_T_102 : _GEN_2809; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2842 = 5'h8 == rd ? _next_reg_T_102 : _GEN_2810; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2843 = 5'h9 == rd ? _next_reg_T_102 : _GEN_2811; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2844 = 5'ha == rd ? _next_reg_T_102 : _GEN_2812; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2845 = 5'hb == rd ? _next_reg_T_102 : _GEN_2813; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2846 = 5'hc == rd ? _next_reg_T_102 : _GEN_2814; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2847 = 5'hd == rd ? _next_reg_T_102 : _GEN_2815; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2848 = 5'he == rd ? _next_reg_T_102 : _GEN_2816; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2849 = 5'hf == rd ? _next_reg_T_102 : _GEN_2817; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2850 = 5'h10 == rd ? _next_reg_T_102 : _GEN_2818; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2851 = 5'h11 == rd ? _next_reg_T_102 : _GEN_2819; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2852 = 5'h12 == rd ? _next_reg_T_102 : _GEN_2820; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2853 = 5'h13 == rd ? _next_reg_T_102 : _GEN_2821; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2854 = 5'h14 == rd ? _next_reg_T_102 : _GEN_2822; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2855 = 5'h15 == rd ? _next_reg_T_102 : _GEN_2823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2856 = 5'h16 == rd ? _next_reg_T_102 : _GEN_2824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2857 = 5'h17 == rd ? _next_reg_T_102 : _GEN_2825; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2858 = 5'h18 == rd ? _next_reg_T_102 : _GEN_2826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2859 = 5'h19 == rd ? _next_reg_T_102 : _GEN_2827; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2860 = 5'h1a == rd ? _next_reg_T_102 : _GEN_2828; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2861 = 5'h1b == rd ? _next_reg_T_102 : _GEN_2829; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2862 = 5'h1c == rd ? _next_reg_T_102 : _GEN_2830; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2863 = 5'h1d == rd ? _next_reg_T_102 : _GEN_2831; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2864 = 5'h1e == rd ? _next_reg_T_102 : _GEN_2832; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2865 = 5'h1f == rd ? _next_reg_T_102 : _GEN_2833; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_2874 = _T_563 ? _GEN_2835 : _GEN_2803; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2875 = _T_563 ? _GEN_2836 : _GEN_2804; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2876 = _T_563 ? _GEN_2837 : _GEN_2805; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2877 = _T_563 ? _GEN_2838 : _GEN_2806; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2878 = _T_563 ? _GEN_2839 : _GEN_2807; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2879 = _T_563 ? _GEN_2840 : _GEN_2808; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2880 = _T_563 ? _GEN_2841 : _GEN_2809; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2881 = _T_563 ? _GEN_2842 : _GEN_2810; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2882 = _T_563 ? _GEN_2843 : _GEN_2811; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2883 = _T_563 ? _GEN_2844 : _GEN_2812; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2884 = _T_563 ? _GEN_2845 : _GEN_2813; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2885 = _T_563 ? _GEN_2846 : _GEN_2814; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2886 = _T_563 ? _GEN_2847 : _GEN_2815; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2887 = _T_563 ? _GEN_2848 : _GEN_2816; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2888 = _T_563 ? _GEN_2849 : _GEN_2817; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2889 = _T_563 ? _GEN_2850 : _GEN_2818; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2890 = _T_563 ? _GEN_2851 : _GEN_2819; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2891 = _T_563 ? _GEN_2852 : _GEN_2820; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2892 = _T_563 ? _GEN_2853 : _GEN_2821; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2893 = _T_563 ? _GEN_2854 : _GEN_2822; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2894 = _T_563 ? _GEN_2855 : _GEN_2823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2895 = _T_563 ? _GEN_2856 : _GEN_2824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2896 = _T_563 ? _GEN_2857 : _GEN_2825; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2897 = _T_563 ? _GEN_2858 : _GEN_2826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2898 = _T_563 ? _GEN_2859 : _GEN_2827; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2899 = _T_563 ? _GEN_2860 : _GEN_2828; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2900 = _T_563 ? _GEN_2861 : _GEN_2829; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2901 = _T_563 ? _GEN_2862 : _GEN_2830; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2902 = _T_563 ? _GEN_2863 : _GEN_2831; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2903 = _T_563 ? _GEN_2864 : _GEN_2832; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_2904 = _T_563 ? _GEN_2865 : _GEN_2833; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [31:0] _next_reg_T_105 = _GEN_31[31:0] >> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:78]
  wire  next_reg_signBit_5 = _next_reg_T_105[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_107 = next_reg_signBit_5 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_108 = {_next_reg_T_107,_next_reg_T_105}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_2906 = 5'h1 == rd ? _next_reg_T_108 : _GEN_2874; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2907 = 5'h2 == rd ? _next_reg_T_108 : _GEN_2875; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2908 = 5'h3 == rd ? _next_reg_T_108 : _GEN_2876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2909 = 5'h4 == rd ? _next_reg_T_108 : _GEN_2877; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2910 = 5'h5 == rd ? _next_reg_T_108 : _GEN_2878; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2911 = 5'h6 == rd ? _next_reg_T_108 : _GEN_2879; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2912 = 5'h7 == rd ? _next_reg_T_108 : _GEN_2880; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2913 = 5'h8 == rd ? _next_reg_T_108 : _GEN_2881; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2914 = 5'h9 == rd ? _next_reg_T_108 : _GEN_2882; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2915 = 5'ha == rd ? _next_reg_T_108 : _GEN_2883; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2916 = 5'hb == rd ? _next_reg_T_108 : _GEN_2884; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2917 = 5'hc == rd ? _next_reg_T_108 : _GEN_2885; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2918 = 5'hd == rd ? _next_reg_T_108 : _GEN_2886; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2919 = 5'he == rd ? _next_reg_T_108 : _GEN_2887; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2920 = 5'hf == rd ? _next_reg_T_108 : _GEN_2888; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2921 = 5'h10 == rd ? _next_reg_T_108 : _GEN_2889; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2922 = 5'h11 == rd ? _next_reg_T_108 : _GEN_2890; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2923 = 5'h12 == rd ? _next_reg_T_108 : _GEN_2891; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2924 = 5'h13 == rd ? _next_reg_T_108 : _GEN_2892; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2925 = 5'h14 == rd ? _next_reg_T_108 : _GEN_2893; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2926 = 5'h15 == rd ? _next_reg_T_108 : _GEN_2894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2927 = 5'h16 == rd ? _next_reg_T_108 : _GEN_2895; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2928 = 5'h17 == rd ? _next_reg_T_108 : _GEN_2896; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2929 = 5'h18 == rd ? _next_reg_T_108 : _GEN_2897; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2930 = 5'h19 == rd ? _next_reg_T_108 : _GEN_2898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2931 = 5'h1a == rd ? _next_reg_T_108 : _GEN_2899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2932 = 5'h1b == rd ? _next_reg_T_108 : _GEN_2900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2933 = 5'h1c == rd ? _next_reg_T_108 : _GEN_2901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2934 = 5'h1d == rd ? _next_reg_T_108 : _GEN_2902; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2935 = 5'h1e == rd ? _next_reg_T_108 : _GEN_2903; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2936 = 5'h1f == rd ? _next_reg_T_108 : _GEN_2904; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_2945 = _T_569 ? _GEN_2906 : _GEN_2874; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2946 = _T_569 ? _GEN_2907 : _GEN_2875; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2947 = _T_569 ? _GEN_2908 : _GEN_2876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2948 = _T_569 ? _GEN_2909 : _GEN_2877; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2949 = _T_569 ? _GEN_2910 : _GEN_2878; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2950 = _T_569 ? _GEN_2911 : _GEN_2879; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2951 = _T_569 ? _GEN_2912 : _GEN_2880; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2952 = _T_569 ? _GEN_2913 : _GEN_2881; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2953 = _T_569 ? _GEN_2914 : _GEN_2882; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2954 = _T_569 ? _GEN_2915 : _GEN_2883; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2955 = _T_569 ? _GEN_2916 : _GEN_2884; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2956 = _T_569 ? _GEN_2917 : _GEN_2885; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2957 = _T_569 ? _GEN_2918 : _GEN_2886; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2958 = _T_569 ? _GEN_2919 : _GEN_2887; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2959 = _T_569 ? _GEN_2920 : _GEN_2888; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2960 = _T_569 ? _GEN_2921 : _GEN_2889; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2961 = _T_569 ? _GEN_2922 : _GEN_2890; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2962 = _T_569 ? _GEN_2923 : _GEN_2891; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2963 = _T_569 ? _GEN_2924 : _GEN_2892; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2964 = _T_569 ? _GEN_2925 : _GEN_2893; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2965 = _T_569 ? _GEN_2926 : _GEN_2894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2966 = _T_569 ? _GEN_2927 : _GEN_2895; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2967 = _T_569 ? _GEN_2928 : _GEN_2896; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2968 = _T_569 ? _GEN_2929 : _GEN_2897; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2969 = _T_569 ? _GEN_2930 : _GEN_2898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2970 = _T_569 ? _GEN_2931 : _GEN_2899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2971 = _T_569 ? _GEN_2932 : _GEN_2900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2972 = _T_569 ? _GEN_2933 : _GEN_2901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2973 = _T_569 ? _GEN_2934 : _GEN_2902; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2974 = _T_569 ? _GEN_2935 : _GEN_2903; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_2975 = _T_569 ? _GEN_2936 : _GEN_2904; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [31:0] _next_reg_T_110 = _GEN_31[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:79]
  wire [31:0] _next_reg_T_113 = $signed(_next_reg_T_110) >>> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:100]
  wire  next_reg_signBit_6 = _next_reg_T_113[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_115 = next_reg_signBit_6 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_116 = {_next_reg_T_115,_next_reg_T_113}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_2977 = 5'h1 == rd ? _next_reg_T_116 : _GEN_2945; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2978 = 5'h2 == rd ? _next_reg_T_116 : _GEN_2946; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2979 = 5'h3 == rd ? _next_reg_T_116 : _GEN_2947; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2980 = 5'h4 == rd ? _next_reg_T_116 : _GEN_2948; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2981 = 5'h5 == rd ? _next_reg_T_116 : _GEN_2949; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2982 = 5'h6 == rd ? _next_reg_T_116 : _GEN_2950; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2983 = 5'h7 == rd ? _next_reg_T_116 : _GEN_2951; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2984 = 5'h8 == rd ? _next_reg_T_116 : _GEN_2952; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2985 = 5'h9 == rd ? _next_reg_T_116 : _GEN_2953; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2986 = 5'ha == rd ? _next_reg_T_116 : _GEN_2954; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2987 = 5'hb == rd ? _next_reg_T_116 : _GEN_2955; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2988 = 5'hc == rd ? _next_reg_T_116 : _GEN_2956; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2989 = 5'hd == rd ? _next_reg_T_116 : _GEN_2957; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2990 = 5'he == rd ? _next_reg_T_116 : _GEN_2958; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2991 = 5'hf == rd ? _next_reg_T_116 : _GEN_2959; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2992 = 5'h10 == rd ? _next_reg_T_116 : _GEN_2960; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2993 = 5'h11 == rd ? _next_reg_T_116 : _GEN_2961; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2994 = 5'h12 == rd ? _next_reg_T_116 : _GEN_2962; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2995 = 5'h13 == rd ? _next_reg_T_116 : _GEN_2963; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2996 = 5'h14 == rd ? _next_reg_T_116 : _GEN_2964; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2997 = 5'h15 == rd ? _next_reg_T_116 : _GEN_2965; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2998 = 5'h16 == rd ? _next_reg_T_116 : _GEN_2966; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_2999 = 5'h17 == rd ? _next_reg_T_116 : _GEN_2967; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_3000 = 5'h18 == rd ? _next_reg_T_116 : _GEN_2968; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_3001 = 5'h19 == rd ? _next_reg_T_116 : _GEN_2969; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_3002 = 5'h1a == rd ? _next_reg_T_116 : _GEN_2970; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_3003 = 5'h1b == rd ? _next_reg_T_116 : _GEN_2971; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_3004 = 5'h1c == rd ? _next_reg_T_116 : _GEN_2972; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_3005 = 5'h1d == rd ? _next_reg_T_116 : _GEN_2973; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_3006 = 5'h1e == rd ? _next_reg_T_116 : _GEN_2974; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_3007 = 5'h1f == rd ? _next_reg_T_116 : _GEN_2975; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_3016 = _T_575 ? _GEN_2977 : _GEN_2945; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3017 = _T_575 ? _GEN_2978 : _GEN_2946; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3018 = _T_575 ? _GEN_2979 : _GEN_2947; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3019 = _T_575 ? _GEN_2980 : _GEN_2948; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3020 = _T_575 ? _GEN_2981 : _GEN_2949; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3021 = _T_575 ? _GEN_2982 : _GEN_2950; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3022 = _T_575 ? _GEN_2983 : _GEN_2951; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3023 = _T_575 ? _GEN_2984 : _GEN_2952; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3024 = _T_575 ? _GEN_2985 : _GEN_2953; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3025 = _T_575 ? _GEN_2986 : _GEN_2954; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3026 = _T_575 ? _GEN_2987 : _GEN_2955; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3027 = _T_575 ? _GEN_2988 : _GEN_2956; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3028 = _T_575 ? _GEN_2989 : _GEN_2957; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3029 = _T_575 ? _GEN_2990 : _GEN_2958; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3030 = _T_575 ? _GEN_2991 : _GEN_2959; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3031 = _T_575 ? _GEN_2992 : _GEN_2960; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3032 = _T_575 ? _GEN_2993 : _GEN_2961; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3033 = _T_575 ? _GEN_2994 : _GEN_2962; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3034 = _T_575 ? _GEN_2995 : _GEN_2963; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3035 = _T_575 ? _GEN_2996 : _GEN_2964; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3036 = _T_575 ? _GEN_2997 : _GEN_2965; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3037 = _T_575 ? _GEN_2998 : _GEN_2966; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3038 = _T_575 ? _GEN_2999 : _GEN_2967; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3039 = _T_575 ? _GEN_3000 : _GEN_2968; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3040 = _T_575 ? _GEN_3001 : _GEN_2969; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3041 = _T_575 ? _GEN_3002 : _GEN_2970; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3042 = _T_575 ? _GEN_3003 : _GEN_2971; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3043 = _T_575 ? _GEN_3004 : _GEN_2972; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3044 = _T_575 ? _GEN_3005 : _GEN_2973; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3045 = _T_575 ? _GEN_3006 : _GEN_2974; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_3046 = _T_575 ? _GEN_3007 : _GEN_2975; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [126:0] _GEN_71 = {{63'd0}, _GEN_31}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:61]
  wire [126:0] _next_reg_T_118 = _GEN_71 << _GEN_840[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:61]
  wire [63:0] _GEN_3048 = 5'h1 == rd ? _next_reg_T_118[63:0] : _GEN_3016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3049 = 5'h2 == rd ? _next_reg_T_118[63:0] : _GEN_3017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3050 = 5'h3 == rd ? _next_reg_T_118[63:0] : _GEN_3018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3051 = 5'h4 == rd ? _next_reg_T_118[63:0] : _GEN_3019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3052 = 5'h5 == rd ? _next_reg_T_118[63:0] : _GEN_3020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3053 = 5'h6 == rd ? _next_reg_T_118[63:0] : _GEN_3021; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3054 = 5'h7 == rd ? _next_reg_T_118[63:0] : _GEN_3022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3055 = 5'h8 == rd ? _next_reg_T_118[63:0] : _GEN_3023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3056 = 5'h9 == rd ? _next_reg_T_118[63:0] : _GEN_3024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3057 = 5'ha == rd ? _next_reg_T_118[63:0] : _GEN_3025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3058 = 5'hb == rd ? _next_reg_T_118[63:0] : _GEN_3026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3059 = 5'hc == rd ? _next_reg_T_118[63:0] : _GEN_3027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3060 = 5'hd == rd ? _next_reg_T_118[63:0] : _GEN_3028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3061 = 5'he == rd ? _next_reg_T_118[63:0] : _GEN_3029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3062 = 5'hf == rd ? _next_reg_T_118[63:0] : _GEN_3030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3063 = 5'h10 == rd ? _next_reg_T_118[63:0] : _GEN_3031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3064 = 5'h11 == rd ? _next_reg_T_118[63:0] : _GEN_3032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3065 = 5'h12 == rd ? _next_reg_T_118[63:0] : _GEN_3033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3066 = 5'h13 == rd ? _next_reg_T_118[63:0] : _GEN_3034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3067 = 5'h14 == rd ? _next_reg_T_118[63:0] : _GEN_3035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3068 = 5'h15 == rd ? _next_reg_T_118[63:0] : _GEN_3036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3069 = 5'h16 == rd ? _next_reg_T_118[63:0] : _GEN_3037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3070 = 5'h17 == rd ? _next_reg_T_118[63:0] : _GEN_3038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3071 = 5'h18 == rd ? _next_reg_T_118[63:0] : _GEN_3039; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3072 = 5'h19 == rd ? _next_reg_T_118[63:0] : _GEN_3040; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3073 = 5'h1a == rd ? _next_reg_T_118[63:0] : _GEN_3041; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3074 = 5'h1b == rd ? _next_reg_T_118[63:0] : _GEN_3042; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3075 = 5'h1c == rd ? _next_reg_T_118[63:0] : _GEN_3043; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3076 = 5'h1d == rd ? _next_reg_T_118[63:0] : _GEN_3044; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3077 = 5'h1e == rd ? _next_reg_T_118[63:0] : _GEN_3045; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3078 = 5'h1f == rd ? _next_reg_T_118[63:0] : _GEN_3046; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_3087 = _T_581 ? _GEN_3048 : _GEN_3016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3088 = _T_581 ? _GEN_3049 : _GEN_3017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3089 = _T_581 ? _GEN_3050 : _GEN_3018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3090 = _T_581 ? _GEN_3051 : _GEN_3019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3091 = _T_581 ? _GEN_3052 : _GEN_3020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3092 = _T_581 ? _GEN_3053 : _GEN_3021; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3093 = _T_581 ? _GEN_3054 : _GEN_3022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3094 = _T_581 ? _GEN_3055 : _GEN_3023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3095 = _T_581 ? _GEN_3056 : _GEN_3024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3096 = _T_581 ? _GEN_3057 : _GEN_3025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3097 = _T_581 ? _GEN_3058 : _GEN_3026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3098 = _T_581 ? _GEN_3059 : _GEN_3027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3099 = _T_581 ? _GEN_3060 : _GEN_3028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3100 = _T_581 ? _GEN_3061 : _GEN_3029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3101 = _T_581 ? _GEN_3062 : _GEN_3030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3102 = _T_581 ? _GEN_3063 : _GEN_3031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3103 = _T_581 ? _GEN_3064 : _GEN_3032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3104 = _T_581 ? _GEN_3065 : _GEN_3033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3105 = _T_581 ? _GEN_3066 : _GEN_3034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3106 = _T_581 ? _GEN_3067 : _GEN_3035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3107 = _T_581 ? _GEN_3068 : _GEN_3036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3108 = _T_581 ? _GEN_3069 : _GEN_3037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3109 = _T_581 ? _GEN_3070 : _GEN_3038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3110 = _T_581 ? _GEN_3071 : _GEN_3039; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3111 = _T_581 ? _GEN_3072 : _GEN_3040; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3112 = _T_581 ? _GEN_3073 : _GEN_3041; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3113 = _T_581 ? _GEN_3074 : _GEN_3042; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3114 = _T_581 ? _GEN_3075 : _GEN_3043; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3115 = _T_581 ? _GEN_3076 : _GEN_3044; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3116 = _T_581 ? _GEN_3077 : _GEN_3045; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_3117 = _T_581 ? _GEN_3078 : _GEN_3046; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _next_reg_T_120 = _GEN_31 >> _GEN_840[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:61]
  wire [63:0] _GEN_3119 = 5'h1 == rd ? _next_reg_T_120 : _GEN_3087; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3120 = 5'h2 == rd ? _next_reg_T_120 : _GEN_3088; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3121 = 5'h3 == rd ? _next_reg_T_120 : _GEN_3089; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3122 = 5'h4 == rd ? _next_reg_T_120 : _GEN_3090; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3123 = 5'h5 == rd ? _next_reg_T_120 : _GEN_3091; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3124 = 5'h6 == rd ? _next_reg_T_120 : _GEN_3092; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3125 = 5'h7 == rd ? _next_reg_T_120 : _GEN_3093; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3126 = 5'h8 == rd ? _next_reg_T_120 : _GEN_3094; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3127 = 5'h9 == rd ? _next_reg_T_120 : _GEN_3095; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3128 = 5'ha == rd ? _next_reg_T_120 : _GEN_3096; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3129 = 5'hb == rd ? _next_reg_T_120 : _GEN_3097; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3130 = 5'hc == rd ? _next_reg_T_120 : _GEN_3098; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3131 = 5'hd == rd ? _next_reg_T_120 : _GEN_3099; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3132 = 5'he == rd ? _next_reg_T_120 : _GEN_3100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3133 = 5'hf == rd ? _next_reg_T_120 : _GEN_3101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3134 = 5'h10 == rd ? _next_reg_T_120 : _GEN_3102; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3135 = 5'h11 == rd ? _next_reg_T_120 : _GEN_3103; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3136 = 5'h12 == rd ? _next_reg_T_120 : _GEN_3104; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3137 = 5'h13 == rd ? _next_reg_T_120 : _GEN_3105; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3138 = 5'h14 == rd ? _next_reg_T_120 : _GEN_3106; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3139 = 5'h15 == rd ? _next_reg_T_120 : _GEN_3107; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3140 = 5'h16 == rd ? _next_reg_T_120 : _GEN_3108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3141 = 5'h17 == rd ? _next_reg_T_120 : _GEN_3109; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3142 = 5'h18 == rd ? _next_reg_T_120 : _GEN_3110; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3143 = 5'h19 == rd ? _next_reg_T_120 : _GEN_3111; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3144 = 5'h1a == rd ? _next_reg_T_120 : _GEN_3112; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3145 = 5'h1b == rd ? _next_reg_T_120 : _GEN_3113; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3146 = 5'h1c == rd ? _next_reg_T_120 : _GEN_3114; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3147 = 5'h1d == rd ? _next_reg_T_120 : _GEN_3115; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3148 = 5'h1e == rd ? _next_reg_T_120 : _GEN_3116; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3149 = 5'h1f == rd ? _next_reg_T_120 : _GEN_3117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_3158 = _T_588 ? _GEN_3119 : _GEN_3087; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3159 = _T_588 ? _GEN_3120 : _GEN_3088; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3160 = _T_588 ? _GEN_3121 : _GEN_3089; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3161 = _T_588 ? _GEN_3122 : _GEN_3090; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3162 = _T_588 ? _GEN_3123 : _GEN_3091; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3163 = _T_588 ? _GEN_3124 : _GEN_3092; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3164 = _T_588 ? _GEN_3125 : _GEN_3093; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3165 = _T_588 ? _GEN_3126 : _GEN_3094; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3166 = _T_588 ? _GEN_3127 : _GEN_3095; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3167 = _T_588 ? _GEN_3128 : _GEN_3096; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3168 = _T_588 ? _GEN_3129 : _GEN_3097; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3169 = _T_588 ? _GEN_3130 : _GEN_3098; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3170 = _T_588 ? _GEN_3131 : _GEN_3099; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3171 = _T_588 ? _GEN_3132 : _GEN_3100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3172 = _T_588 ? _GEN_3133 : _GEN_3101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3173 = _T_588 ? _GEN_3134 : _GEN_3102; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3174 = _T_588 ? _GEN_3135 : _GEN_3103; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3175 = _T_588 ? _GEN_3136 : _GEN_3104; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3176 = _T_588 ? _GEN_3137 : _GEN_3105; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3177 = _T_588 ? _GEN_3138 : _GEN_3106; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3178 = _T_588 ? _GEN_3139 : _GEN_3107; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3179 = _T_588 ? _GEN_3140 : _GEN_3108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3180 = _T_588 ? _GEN_3141 : _GEN_3109; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3181 = _T_588 ? _GEN_3142 : _GEN_3110; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3182 = _T_588 ? _GEN_3143 : _GEN_3111; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3183 = _T_588 ? _GEN_3144 : _GEN_3112; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3184 = _T_588 ? _GEN_3145 : _GEN_3113; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3185 = _T_588 ? _GEN_3146 : _GEN_3114; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3186 = _T_588 ? _GEN_3147 : _GEN_3115; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3187 = _T_588 ? _GEN_3148 : _GEN_3116; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_3188 = _T_588 ? _GEN_3149 : _GEN_3117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _next_reg_T_124 = $signed(_T_300) >>> _GEN_840[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:92]
  wire [63:0] _GEN_3190 = 5'h1 == rd ? _next_reg_T_124 : _GEN_3158; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3191 = 5'h2 == rd ? _next_reg_T_124 : _GEN_3159; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3192 = 5'h3 == rd ? _next_reg_T_124 : _GEN_3160; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3193 = 5'h4 == rd ? _next_reg_T_124 : _GEN_3161; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3194 = 5'h5 == rd ? _next_reg_T_124 : _GEN_3162; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3195 = 5'h6 == rd ? _next_reg_T_124 : _GEN_3163; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3196 = 5'h7 == rd ? _next_reg_T_124 : _GEN_3164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3197 = 5'h8 == rd ? _next_reg_T_124 : _GEN_3165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3198 = 5'h9 == rd ? _next_reg_T_124 : _GEN_3166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3199 = 5'ha == rd ? _next_reg_T_124 : _GEN_3167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3200 = 5'hb == rd ? _next_reg_T_124 : _GEN_3168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3201 = 5'hc == rd ? _next_reg_T_124 : _GEN_3169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3202 = 5'hd == rd ? _next_reg_T_124 : _GEN_3170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3203 = 5'he == rd ? _next_reg_T_124 : _GEN_3171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3204 = 5'hf == rd ? _next_reg_T_124 : _GEN_3172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3205 = 5'h10 == rd ? _next_reg_T_124 : _GEN_3173; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3206 = 5'h11 == rd ? _next_reg_T_124 : _GEN_3174; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3207 = 5'h12 == rd ? _next_reg_T_124 : _GEN_3175; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3208 = 5'h13 == rd ? _next_reg_T_124 : _GEN_3176; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3209 = 5'h14 == rd ? _next_reg_T_124 : _GEN_3177; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3210 = 5'h15 == rd ? _next_reg_T_124 : _GEN_3178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3211 = 5'h16 == rd ? _next_reg_T_124 : _GEN_3179; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3212 = 5'h17 == rd ? _next_reg_T_124 : _GEN_3180; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3213 = 5'h18 == rd ? _next_reg_T_124 : _GEN_3181; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3214 = 5'h19 == rd ? _next_reg_T_124 : _GEN_3182; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3215 = 5'h1a == rd ? _next_reg_T_124 : _GEN_3183; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3216 = 5'h1b == rd ? _next_reg_T_124 : _GEN_3184; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3217 = 5'h1c == rd ? _next_reg_T_124 : _GEN_3185; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3218 = 5'h1d == rd ? _next_reg_T_124 : _GEN_3186; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3219 = 5'h1e == rd ? _next_reg_T_124 : _GEN_3187; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3220 = 5'h1f == rd ? _next_reg_T_124 : _GEN_3188; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_3229 = _T_595 ? _GEN_3190 : _GEN_3158; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3230 = _T_595 ? _GEN_3191 : _GEN_3159; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3231 = _T_595 ? _GEN_3192 : _GEN_3160; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3232 = _T_595 ? _GEN_3193 : _GEN_3161; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3233 = _T_595 ? _GEN_3194 : _GEN_3162; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3234 = _T_595 ? _GEN_3195 : _GEN_3163; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3235 = _T_595 ? _GEN_3196 : _GEN_3164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3236 = _T_595 ? _GEN_3197 : _GEN_3165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3237 = _T_595 ? _GEN_3198 : _GEN_3166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3238 = _T_595 ? _GEN_3199 : _GEN_3167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3239 = _T_595 ? _GEN_3200 : _GEN_3168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3240 = _T_595 ? _GEN_3201 : _GEN_3169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3241 = _T_595 ? _GEN_3202 : _GEN_3170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3242 = _T_595 ? _GEN_3203 : _GEN_3171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3243 = _T_595 ? _GEN_3204 : _GEN_3172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3244 = _T_595 ? _GEN_3205 : _GEN_3173; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3245 = _T_595 ? _GEN_3206 : _GEN_3174; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3246 = _T_595 ? _GEN_3207 : _GEN_3175; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3247 = _T_595 ? _GEN_3208 : _GEN_3176; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3248 = _T_595 ? _GEN_3209 : _GEN_3177; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3249 = _T_595 ? _GEN_3210 : _GEN_3178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3250 = _T_595 ? _GEN_3211 : _GEN_3179; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3251 = _T_595 ? _GEN_3212 : _GEN_3180; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3252 = _T_595 ? _GEN_3213 : _GEN_3181; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3253 = _T_595 ? _GEN_3214 : _GEN_3182; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3254 = _T_595 ? _GEN_3215 : _GEN_3183; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3255 = _T_595 ? _GEN_3216 : _GEN_3184; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3256 = _T_595 ? _GEN_3217 : _GEN_3185; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3257 = _T_595 ? _GEN_3218 : _GEN_3186; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3258 = _T_595 ? _GEN_3219 : _GEN_3187; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_3259 = _T_595 ? _GEN_3220 : _GEN_3188; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [31:0] _next_reg_T_128 = _GEN_31[31:0] + _GEN_840[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:78]
  wire  next_reg_signBit_7 = _next_reg_T_128[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_131 = next_reg_signBit_7 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_132 = {_next_reg_T_131,_next_reg_T_128}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_3261 = 5'h1 == rd ? _next_reg_T_132 : _GEN_3229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3262 = 5'h2 == rd ? _next_reg_T_132 : _GEN_3230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3263 = 5'h3 == rd ? _next_reg_T_132 : _GEN_3231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3264 = 5'h4 == rd ? _next_reg_T_132 : _GEN_3232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3265 = 5'h5 == rd ? _next_reg_T_132 : _GEN_3233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3266 = 5'h6 == rd ? _next_reg_T_132 : _GEN_3234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3267 = 5'h7 == rd ? _next_reg_T_132 : _GEN_3235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3268 = 5'h8 == rd ? _next_reg_T_132 : _GEN_3236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3269 = 5'h9 == rd ? _next_reg_T_132 : _GEN_3237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3270 = 5'ha == rd ? _next_reg_T_132 : _GEN_3238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3271 = 5'hb == rd ? _next_reg_T_132 : _GEN_3239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3272 = 5'hc == rd ? _next_reg_T_132 : _GEN_3240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3273 = 5'hd == rd ? _next_reg_T_132 : _GEN_3241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3274 = 5'he == rd ? _next_reg_T_132 : _GEN_3242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3275 = 5'hf == rd ? _next_reg_T_132 : _GEN_3243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3276 = 5'h10 == rd ? _next_reg_T_132 : _GEN_3244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3277 = 5'h11 == rd ? _next_reg_T_132 : _GEN_3245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3278 = 5'h12 == rd ? _next_reg_T_132 : _GEN_3246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3279 = 5'h13 == rd ? _next_reg_T_132 : _GEN_3247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3280 = 5'h14 == rd ? _next_reg_T_132 : _GEN_3248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3281 = 5'h15 == rd ? _next_reg_T_132 : _GEN_3249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3282 = 5'h16 == rd ? _next_reg_T_132 : _GEN_3250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3283 = 5'h17 == rd ? _next_reg_T_132 : _GEN_3251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3284 = 5'h18 == rd ? _next_reg_T_132 : _GEN_3252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3285 = 5'h19 == rd ? _next_reg_T_132 : _GEN_3253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3286 = 5'h1a == rd ? _next_reg_T_132 : _GEN_3254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3287 = 5'h1b == rd ? _next_reg_T_132 : _GEN_3255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3288 = 5'h1c == rd ? _next_reg_T_132 : _GEN_3256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3289 = 5'h1d == rd ? _next_reg_T_132 : _GEN_3257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3290 = 5'h1e == rd ? _next_reg_T_132 : _GEN_3258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3291 = 5'h1f == rd ? _next_reg_T_132 : _GEN_3259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_3300 = _T_602 ? _GEN_3261 : _GEN_3229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3301 = _T_602 ? _GEN_3262 : _GEN_3230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3302 = _T_602 ? _GEN_3263 : _GEN_3231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3303 = _T_602 ? _GEN_3264 : _GEN_3232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3304 = _T_602 ? _GEN_3265 : _GEN_3233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3305 = _T_602 ? _GEN_3266 : _GEN_3234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3306 = _T_602 ? _GEN_3267 : _GEN_3235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3307 = _T_602 ? _GEN_3268 : _GEN_3236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3308 = _T_602 ? _GEN_3269 : _GEN_3237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3309 = _T_602 ? _GEN_3270 : _GEN_3238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3310 = _T_602 ? _GEN_3271 : _GEN_3239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3311 = _T_602 ? _GEN_3272 : _GEN_3240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3312 = _T_602 ? _GEN_3273 : _GEN_3241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3313 = _T_602 ? _GEN_3274 : _GEN_3242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3314 = _T_602 ? _GEN_3275 : _GEN_3243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3315 = _T_602 ? _GEN_3276 : _GEN_3244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3316 = _T_602 ? _GEN_3277 : _GEN_3245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3317 = _T_602 ? _GEN_3278 : _GEN_3246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3318 = _T_602 ? _GEN_3279 : _GEN_3247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3319 = _T_602 ? _GEN_3280 : _GEN_3248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3320 = _T_602 ? _GEN_3281 : _GEN_3249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3321 = _T_602 ? _GEN_3282 : _GEN_3250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3322 = _T_602 ? _GEN_3283 : _GEN_3251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3323 = _T_602 ? _GEN_3284 : _GEN_3252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3324 = _T_602 ? _GEN_3285 : _GEN_3253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3325 = _T_602 ? _GEN_3286 : _GEN_3254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3326 = _T_602 ? _GEN_3287 : _GEN_3255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3327 = _T_602 ? _GEN_3288 : _GEN_3256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3328 = _T_602 ? _GEN_3289 : _GEN_3257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3329 = _T_602 ? _GEN_3290 : _GEN_3258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_3330 = _T_602 ? _GEN_3291 : _GEN_3259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [62:0] _GEN_103 = {{31'd0}, _GEN_31[31:0]}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:78]
  wire [62:0] _next_reg_T_135 = _GEN_103 << _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:78]
  wire  next_reg_signBit_8 = _next_reg_T_135[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_138 = next_reg_signBit_8 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_139 = {_next_reg_T_138,_next_reg_T_135[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_3332 = 5'h1 == rd ? _next_reg_T_139 : _GEN_3300; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3333 = 5'h2 == rd ? _next_reg_T_139 : _GEN_3301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3334 = 5'h3 == rd ? _next_reg_T_139 : _GEN_3302; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3335 = 5'h4 == rd ? _next_reg_T_139 : _GEN_3303; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3336 = 5'h5 == rd ? _next_reg_T_139 : _GEN_3304; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3337 = 5'h6 == rd ? _next_reg_T_139 : _GEN_3305; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3338 = 5'h7 == rd ? _next_reg_T_139 : _GEN_3306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3339 = 5'h8 == rd ? _next_reg_T_139 : _GEN_3307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3340 = 5'h9 == rd ? _next_reg_T_139 : _GEN_3308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3341 = 5'ha == rd ? _next_reg_T_139 : _GEN_3309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3342 = 5'hb == rd ? _next_reg_T_139 : _GEN_3310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3343 = 5'hc == rd ? _next_reg_T_139 : _GEN_3311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3344 = 5'hd == rd ? _next_reg_T_139 : _GEN_3312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3345 = 5'he == rd ? _next_reg_T_139 : _GEN_3313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3346 = 5'hf == rd ? _next_reg_T_139 : _GEN_3314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3347 = 5'h10 == rd ? _next_reg_T_139 : _GEN_3315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3348 = 5'h11 == rd ? _next_reg_T_139 : _GEN_3316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3349 = 5'h12 == rd ? _next_reg_T_139 : _GEN_3317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3350 = 5'h13 == rd ? _next_reg_T_139 : _GEN_3318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3351 = 5'h14 == rd ? _next_reg_T_139 : _GEN_3319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3352 = 5'h15 == rd ? _next_reg_T_139 : _GEN_3320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3353 = 5'h16 == rd ? _next_reg_T_139 : _GEN_3321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3354 = 5'h17 == rd ? _next_reg_T_139 : _GEN_3322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3355 = 5'h18 == rd ? _next_reg_T_139 : _GEN_3323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3356 = 5'h19 == rd ? _next_reg_T_139 : _GEN_3324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3357 = 5'h1a == rd ? _next_reg_T_139 : _GEN_3325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3358 = 5'h1b == rd ? _next_reg_T_139 : _GEN_3326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3359 = 5'h1c == rd ? _next_reg_T_139 : _GEN_3327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3360 = 5'h1d == rd ? _next_reg_T_139 : _GEN_3328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3361 = 5'h1e == rd ? _next_reg_T_139 : _GEN_3329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3362 = 5'h1f == rd ? _next_reg_T_139 : _GEN_3330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_3371 = _T_609 ? _GEN_3332 : _GEN_3300; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3372 = _T_609 ? _GEN_3333 : _GEN_3301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3373 = _T_609 ? _GEN_3334 : _GEN_3302; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3374 = _T_609 ? _GEN_3335 : _GEN_3303; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3375 = _T_609 ? _GEN_3336 : _GEN_3304; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3376 = _T_609 ? _GEN_3337 : _GEN_3305; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3377 = _T_609 ? _GEN_3338 : _GEN_3306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3378 = _T_609 ? _GEN_3339 : _GEN_3307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3379 = _T_609 ? _GEN_3340 : _GEN_3308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3380 = _T_609 ? _GEN_3341 : _GEN_3309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3381 = _T_609 ? _GEN_3342 : _GEN_3310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3382 = _T_609 ? _GEN_3343 : _GEN_3311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3383 = _T_609 ? _GEN_3344 : _GEN_3312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3384 = _T_609 ? _GEN_3345 : _GEN_3313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3385 = _T_609 ? _GEN_3346 : _GEN_3314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3386 = _T_609 ? _GEN_3347 : _GEN_3315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3387 = _T_609 ? _GEN_3348 : _GEN_3316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3388 = _T_609 ? _GEN_3349 : _GEN_3317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3389 = _T_609 ? _GEN_3350 : _GEN_3318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3390 = _T_609 ? _GEN_3351 : _GEN_3319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3391 = _T_609 ? _GEN_3352 : _GEN_3320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3392 = _T_609 ? _GEN_3353 : _GEN_3321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3393 = _T_609 ? _GEN_3354 : _GEN_3322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3394 = _T_609 ? _GEN_3355 : _GEN_3323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3395 = _T_609 ? _GEN_3356 : _GEN_3324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3396 = _T_609 ? _GEN_3357 : _GEN_3325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3397 = _T_609 ? _GEN_3358 : _GEN_3326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3398 = _T_609 ? _GEN_3359 : _GEN_3327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3399 = _T_609 ? _GEN_3360 : _GEN_3328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3400 = _T_609 ? _GEN_3361 : _GEN_3329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_3401 = _T_609 ? _GEN_3362 : _GEN_3330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [31:0] _next_reg_T_142 = _GEN_31[31:0] >> _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:78]
  wire  next_reg_signBit_9 = _next_reg_T_142[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_145 = next_reg_signBit_9 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_146 = {_next_reg_T_145,_next_reg_T_142}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_3403 = 5'h1 == rd ? _next_reg_T_146 : _GEN_3371; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3404 = 5'h2 == rd ? _next_reg_T_146 : _GEN_3372; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3405 = 5'h3 == rd ? _next_reg_T_146 : _GEN_3373; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3406 = 5'h4 == rd ? _next_reg_T_146 : _GEN_3374; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3407 = 5'h5 == rd ? _next_reg_T_146 : _GEN_3375; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3408 = 5'h6 == rd ? _next_reg_T_146 : _GEN_3376; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3409 = 5'h7 == rd ? _next_reg_T_146 : _GEN_3377; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3410 = 5'h8 == rd ? _next_reg_T_146 : _GEN_3378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3411 = 5'h9 == rd ? _next_reg_T_146 : _GEN_3379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3412 = 5'ha == rd ? _next_reg_T_146 : _GEN_3380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3413 = 5'hb == rd ? _next_reg_T_146 : _GEN_3381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3414 = 5'hc == rd ? _next_reg_T_146 : _GEN_3382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3415 = 5'hd == rd ? _next_reg_T_146 : _GEN_3383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3416 = 5'he == rd ? _next_reg_T_146 : _GEN_3384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3417 = 5'hf == rd ? _next_reg_T_146 : _GEN_3385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3418 = 5'h10 == rd ? _next_reg_T_146 : _GEN_3386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3419 = 5'h11 == rd ? _next_reg_T_146 : _GEN_3387; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3420 = 5'h12 == rd ? _next_reg_T_146 : _GEN_3388; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3421 = 5'h13 == rd ? _next_reg_T_146 : _GEN_3389; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3422 = 5'h14 == rd ? _next_reg_T_146 : _GEN_3390; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3423 = 5'h15 == rd ? _next_reg_T_146 : _GEN_3391; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3424 = 5'h16 == rd ? _next_reg_T_146 : _GEN_3392; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3425 = 5'h17 == rd ? _next_reg_T_146 : _GEN_3393; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3426 = 5'h18 == rd ? _next_reg_T_146 : _GEN_3394; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3427 = 5'h19 == rd ? _next_reg_T_146 : _GEN_3395; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3428 = 5'h1a == rd ? _next_reg_T_146 : _GEN_3396; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3429 = 5'h1b == rd ? _next_reg_T_146 : _GEN_3397; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3430 = 5'h1c == rd ? _next_reg_T_146 : _GEN_3398; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3431 = 5'h1d == rd ? _next_reg_T_146 : _GEN_3399; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3432 = 5'h1e == rd ? _next_reg_T_146 : _GEN_3400; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3433 = 5'h1f == rd ? _next_reg_T_146 : _GEN_3401; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_3442 = _T_616 ? _GEN_3403 : _GEN_3371; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3443 = _T_616 ? _GEN_3404 : _GEN_3372; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3444 = _T_616 ? _GEN_3405 : _GEN_3373; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3445 = _T_616 ? _GEN_3406 : _GEN_3374; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3446 = _T_616 ? _GEN_3407 : _GEN_3375; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3447 = _T_616 ? _GEN_3408 : _GEN_3376; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3448 = _T_616 ? _GEN_3409 : _GEN_3377; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3449 = _T_616 ? _GEN_3410 : _GEN_3378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3450 = _T_616 ? _GEN_3411 : _GEN_3379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3451 = _T_616 ? _GEN_3412 : _GEN_3380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3452 = _T_616 ? _GEN_3413 : _GEN_3381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3453 = _T_616 ? _GEN_3414 : _GEN_3382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3454 = _T_616 ? _GEN_3415 : _GEN_3383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3455 = _T_616 ? _GEN_3416 : _GEN_3384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3456 = _T_616 ? _GEN_3417 : _GEN_3385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3457 = _T_616 ? _GEN_3418 : _GEN_3386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3458 = _T_616 ? _GEN_3419 : _GEN_3387; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3459 = _T_616 ? _GEN_3420 : _GEN_3388; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3460 = _T_616 ? _GEN_3421 : _GEN_3389; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3461 = _T_616 ? _GEN_3422 : _GEN_3390; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3462 = _T_616 ? _GEN_3423 : _GEN_3391; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3463 = _T_616 ? _GEN_3424 : _GEN_3392; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3464 = _T_616 ? _GEN_3425 : _GEN_3393; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3465 = _T_616 ? _GEN_3426 : _GEN_3394; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3466 = _T_616 ? _GEN_3427 : _GEN_3395; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3467 = _T_616 ? _GEN_3428 : _GEN_3396; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3468 = _T_616 ? _GEN_3429 : _GEN_3397; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3469 = _T_616 ? _GEN_3430 : _GEN_3398; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3470 = _T_616 ? _GEN_3431 : _GEN_3399; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3471 = _T_616 ? _GEN_3432 : _GEN_3400; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_3472 = _T_616 ? _GEN_3433 : _GEN_3401; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [31:0] _next_reg_T_150 = _GEN_31[31:0] - _GEN_840[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:78]
  wire  next_reg_signBit_10 = _next_reg_T_150[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_153 = next_reg_signBit_10 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_154 = {_next_reg_T_153,_next_reg_T_150}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_3474 = 5'h1 == rd ? _next_reg_T_154 : _GEN_3442; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3475 = 5'h2 == rd ? _next_reg_T_154 : _GEN_3443; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3476 = 5'h3 == rd ? _next_reg_T_154 : _GEN_3444; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3477 = 5'h4 == rd ? _next_reg_T_154 : _GEN_3445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3478 = 5'h5 == rd ? _next_reg_T_154 : _GEN_3446; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3479 = 5'h6 == rd ? _next_reg_T_154 : _GEN_3447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3480 = 5'h7 == rd ? _next_reg_T_154 : _GEN_3448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3481 = 5'h8 == rd ? _next_reg_T_154 : _GEN_3449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3482 = 5'h9 == rd ? _next_reg_T_154 : _GEN_3450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3483 = 5'ha == rd ? _next_reg_T_154 : _GEN_3451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3484 = 5'hb == rd ? _next_reg_T_154 : _GEN_3452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3485 = 5'hc == rd ? _next_reg_T_154 : _GEN_3453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3486 = 5'hd == rd ? _next_reg_T_154 : _GEN_3454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3487 = 5'he == rd ? _next_reg_T_154 : _GEN_3455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3488 = 5'hf == rd ? _next_reg_T_154 : _GEN_3456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3489 = 5'h10 == rd ? _next_reg_T_154 : _GEN_3457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3490 = 5'h11 == rd ? _next_reg_T_154 : _GEN_3458; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3491 = 5'h12 == rd ? _next_reg_T_154 : _GEN_3459; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3492 = 5'h13 == rd ? _next_reg_T_154 : _GEN_3460; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3493 = 5'h14 == rd ? _next_reg_T_154 : _GEN_3461; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3494 = 5'h15 == rd ? _next_reg_T_154 : _GEN_3462; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3495 = 5'h16 == rd ? _next_reg_T_154 : _GEN_3463; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3496 = 5'h17 == rd ? _next_reg_T_154 : _GEN_3464; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3497 = 5'h18 == rd ? _next_reg_T_154 : _GEN_3465; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3498 = 5'h19 == rd ? _next_reg_T_154 : _GEN_3466; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3499 = 5'h1a == rd ? _next_reg_T_154 : _GEN_3467; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3500 = 5'h1b == rd ? _next_reg_T_154 : _GEN_3468; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3501 = 5'h1c == rd ? _next_reg_T_154 : _GEN_3469; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3502 = 5'h1d == rd ? _next_reg_T_154 : _GEN_3470; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3503 = 5'h1e == rd ? _next_reg_T_154 : _GEN_3471; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3504 = 5'h1f == rd ? _next_reg_T_154 : _GEN_3472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_3513 = _T_623 ? _GEN_3474 : _GEN_3442; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3514 = _T_623 ? _GEN_3475 : _GEN_3443; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3515 = _T_623 ? _GEN_3476 : _GEN_3444; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3516 = _T_623 ? _GEN_3477 : _GEN_3445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3517 = _T_623 ? _GEN_3478 : _GEN_3446; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3518 = _T_623 ? _GEN_3479 : _GEN_3447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3519 = _T_623 ? _GEN_3480 : _GEN_3448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3520 = _T_623 ? _GEN_3481 : _GEN_3449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3521 = _T_623 ? _GEN_3482 : _GEN_3450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3522 = _T_623 ? _GEN_3483 : _GEN_3451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3523 = _T_623 ? _GEN_3484 : _GEN_3452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3524 = _T_623 ? _GEN_3485 : _GEN_3453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3525 = _T_623 ? _GEN_3486 : _GEN_3454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3526 = _T_623 ? _GEN_3487 : _GEN_3455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3527 = _T_623 ? _GEN_3488 : _GEN_3456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3528 = _T_623 ? _GEN_3489 : _GEN_3457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3529 = _T_623 ? _GEN_3490 : _GEN_3458; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3530 = _T_623 ? _GEN_3491 : _GEN_3459; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3531 = _T_623 ? _GEN_3492 : _GEN_3460; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3532 = _T_623 ? _GEN_3493 : _GEN_3461; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3533 = _T_623 ? _GEN_3494 : _GEN_3462; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3534 = _T_623 ? _GEN_3495 : _GEN_3463; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3535 = _T_623 ? _GEN_3496 : _GEN_3464; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3536 = _T_623 ? _GEN_3497 : _GEN_3465; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3537 = _T_623 ? _GEN_3498 : _GEN_3466; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3538 = _T_623 ? _GEN_3499 : _GEN_3467; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3539 = _T_623 ? _GEN_3500 : _GEN_3468; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3540 = _T_623 ? _GEN_3501 : _GEN_3469; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3541 = _T_623 ? _GEN_3502 : _GEN_3470; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3542 = _T_623 ? _GEN_3503 : _GEN_3471; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_3543 = _T_623 ? _GEN_3504 : _GEN_3472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [31:0] _next_reg_T_159 = $signed(_next_reg_T_110) >>> _GEN_840[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:108]
  wire  next_reg_signBit_11 = _next_reg_T_159[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_161 = next_reg_signBit_11 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_162 = {_next_reg_T_161,_next_reg_T_159}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_3545 = 5'h1 == rd ? _next_reg_T_162 : _GEN_3513; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3546 = 5'h2 == rd ? _next_reg_T_162 : _GEN_3514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3547 = 5'h3 == rd ? _next_reg_T_162 : _GEN_3515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3548 = 5'h4 == rd ? _next_reg_T_162 : _GEN_3516; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3549 = 5'h5 == rd ? _next_reg_T_162 : _GEN_3517; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3550 = 5'h6 == rd ? _next_reg_T_162 : _GEN_3518; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3551 = 5'h7 == rd ? _next_reg_T_162 : _GEN_3519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3552 = 5'h8 == rd ? _next_reg_T_162 : _GEN_3520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3553 = 5'h9 == rd ? _next_reg_T_162 : _GEN_3521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3554 = 5'ha == rd ? _next_reg_T_162 : _GEN_3522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3555 = 5'hb == rd ? _next_reg_T_162 : _GEN_3523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3556 = 5'hc == rd ? _next_reg_T_162 : _GEN_3524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3557 = 5'hd == rd ? _next_reg_T_162 : _GEN_3525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3558 = 5'he == rd ? _next_reg_T_162 : _GEN_3526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3559 = 5'hf == rd ? _next_reg_T_162 : _GEN_3527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3560 = 5'h10 == rd ? _next_reg_T_162 : _GEN_3528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3561 = 5'h11 == rd ? _next_reg_T_162 : _GEN_3529; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3562 = 5'h12 == rd ? _next_reg_T_162 : _GEN_3530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3563 = 5'h13 == rd ? _next_reg_T_162 : _GEN_3531; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3564 = 5'h14 == rd ? _next_reg_T_162 : _GEN_3532; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3565 = 5'h15 == rd ? _next_reg_T_162 : _GEN_3533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3566 = 5'h16 == rd ? _next_reg_T_162 : _GEN_3534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3567 = 5'h17 == rd ? _next_reg_T_162 : _GEN_3535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3568 = 5'h18 == rd ? _next_reg_T_162 : _GEN_3536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3569 = 5'h19 == rd ? _next_reg_T_162 : _GEN_3537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3570 = 5'h1a == rd ? _next_reg_T_162 : _GEN_3538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3571 = 5'h1b == rd ? _next_reg_T_162 : _GEN_3539; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3572 = 5'h1c == rd ? _next_reg_T_162 : _GEN_3540; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3573 = 5'h1d == rd ? _next_reg_T_162 : _GEN_3541; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3574 = 5'h1e == rd ? _next_reg_T_162 : _GEN_3542; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3575 = 5'h1f == rd ? _next_reg_T_162 : _GEN_3543; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_3584 = _T_630 ? _GEN_3545 : _GEN_3513; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3585 = _T_630 ? _GEN_3546 : _GEN_3514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3586 = _T_630 ? _GEN_3547 : _GEN_3515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3587 = _T_630 ? _GEN_3548 : _GEN_3516; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3588 = _T_630 ? _GEN_3549 : _GEN_3517; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3589 = _T_630 ? _GEN_3550 : _GEN_3518; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3590 = _T_630 ? _GEN_3551 : _GEN_3519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3591 = _T_630 ? _GEN_3552 : _GEN_3520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3592 = _T_630 ? _GEN_3553 : _GEN_3521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3593 = _T_630 ? _GEN_3554 : _GEN_3522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3594 = _T_630 ? _GEN_3555 : _GEN_3523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3595 = _T_630 ? _GEN_3556 : _GEN_3524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3596 = _T_630 ? _GEN_3557 : _GEN_3525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3597 = _T_630 ? _GEN_3558 : _GEN_3526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3598 = _T_630 ? _GEN_3559 : _GEN_3527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3599 = _T_630 ? _GEN_3560 : _GEN_3528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3600 = _T_630 ? _GEN_3561 : _GEN_3529; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3601 = _T_630 ? _GEN_3562 : _GEN_3530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3602 = _T_630 ? _GEN_3563 : _GEN_3531; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3603 = _T_630 ? _GEN_3564 : _GEN_3532; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3604 = _T_630 ? _GEN_3565 : _GEN_3533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3605 = _T_630 ? _GEN_3566 : _GEN_3534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3606 = _T_630 ? _GEN_3567 : _GEN_3535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3607 = _T_630 ? _GEN_3568 : _GEN_3536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3608 = _T_630 ? _GEN_3569 : _GEN_3537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3609 = _T_630 ? _GEN_3570 : _GEN_3538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3610 = _T_630 ? _GEN_3571 : _GEN_3539; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3611 = _T_630 ? _GEN_3572 : _GEN_3540; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3612 = _T_630 ? _GEN_3573 : _GEN_3541; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3613 = _T_630 ? _GEN_3574 : _GEN_3542; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_3614 = _T_630 ? _GEN_3575 : _GEN_3543; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _next_reg_T_168 = {32'h0,_next_reg_T_65[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [63:0] _GEN_3616 = 5'h1 == rd ? _next_reg_T_168 : _GEN_3584; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3617 = 5'h2 == rd ? _next_reg_T_168 : _GEN_3585; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3618 = 5'h3 == rd ? _next_reg_T_168 : _GEN_3586; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3619 = 5'h4 == rd ? _next_reg_T_168 : _GEN_3587; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3620 = 5'h5 == rd ? _next_reg_T_168 : _GEN_3588; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3621 = 5'h6 == rd ? _next_reg_T_168 : _GEN_3589; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3622 = 5'h7 == rd ? _next_reg_T_168 : _GEN_3590; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3623 = 5'h8 == rd ? _next_reg_T_168 : _GEN_3591; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3624 = 5'h9 == rd ? _next_reg_T_168 : _GEN_3592; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3625 = 5'ha == rd ? _next_reg_T_168 : _GEN_3593; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3626 = 5'hb == rd ? _next_reg_T_168 : _GEN_3594; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3627 = 5'hc == rd ? _next_reg_T_168 : _GEN_3595; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3628 = 5'hd == rd ? _next_reg_T_168 : _GEN_3596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3629 = 5'he == rd ? _next_reg_T_168 : _GEN_3597; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3630 = 5'hf == rd ? _next_reg_T_168 : _GEN_3598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3631 = 5'h10 == rd ? _next_reg_T_168 : _GEN_3599; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3632 = 5'h11 == rd ? _next_reg_T_168 : _GEN_3600; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3633 = 5'h12 == rd ? _next_reg_T_168 : _GEN_3601; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3634 = 5'h13 == rd ? _next_reg_T_168 : _GEN_3602; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3635 = 5'h14 == rd ? _next_reg_T_168 : _GEN_3603; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3636 = 5'h15 == rd ? _next_reg_T_168 : _GEN_3604; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3637 = 5'h16 == rd ? _next_reg_T_168 : _GEN_3605; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3638 = 5'h17 == rd ? _next_reg_T_168 : _GEN_3606; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3639 = 5'h18 == rd ? _next_reg_T_168 : _GEN_3607; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3640 = 5'h19 == rd ? _next_reg_T_168 : _GEN_3608; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3641 = 5'h1a == rd ? _next_reg_T_168 : _GEN_3609; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3642 = 5'h1b == rd ? _next_reg_T_168 : _GEN_3610; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3643 = 5'h1c == rd ? _next_reg_T_168 : _GEN_3611; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3644 = 5'h1d == rd ? _next_reg_T_168 : _GEN_3612; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3645 = 5'h1e == rd ? _next_reg_T_168 : _GEN_3613; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_3646 = 5'h1f == rd ? _next_reg_T_168 : _GEN_3614; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire  _GEN_3647 = _T_667 | _GEN_2421; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [6:0] _GEN_3649 = _T_667 ? 7'h20 : _GEN_2423; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [63:0] _GEN_3651 = _T_667 ? _GEN_3616 : _GEN_3584; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3652 = _T_667 ? _GEN_3617 : _GEN_3585; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3653 = _T_667 ? _GEN_3618 : _GEN_3586; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3654 = _T_667 ? _GEN_3619 : _GEN_3587; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3655 = _T_667 ? _GEN_3620 : _GEN_3588; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3656 = _T_667 ? _GEN_3621 : _GEN_3589; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3657 = _T_667 ? _GEN_3622 : _GEN_3590; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3658 = _T_667 ? _GEN_3623 : _GEN_3591; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3659 = _T_667 ? _GEN_3624 : _GEN_3592; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3660 = _T_667 ? _GEN_3625 : _GEN_3593; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3661 = _T_667 ? _GEN_3626 : _GEN_3594; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3662 = _T_667 ? _GEN_3627 : _GEN_3595; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3663 = _T_667 ? _GEN_3628 : _GEN_3596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3664 = _T_667 ? _GEN_3629 : _GEN_3597; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3665 = _T_667 ? _GEN_3630 : _GEN_3598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3666 = _T_667 ? _GEN_3631 : _GEN_3599; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3667 = _T_667 ? _GEN_3632 : _GEN_3600; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3668 = _T_667 ? _GEN_3633 : _GEN_3601; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3669 = _T_667 ? _GEN_3634 : _GEN_3602; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3670 = _T_667 ? _GEN_3635 : _GEN_3603; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3671 = _T_667 ? _GEN_3636 : _GEN_3604; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3672 = _T_667 ? _GEN_3637 : _GEN_3605; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3673 = _T_667 ? _GEN_3638 : _GEN_3606; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3674 = _T_667 ? _GEN_3639 : _GEN_3607; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3675 = _T_667 ? _GEN_3640 : _GEN_3608; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3676 = _T_667 ? _GEN_3641 : _GEN_3609; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3677 = _T_667 ? _GEN_3642 : _GEN_3610; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3678 = _T_667 ? _GEN_3643 : _GEN_3611; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3679 = _T_667 ? _GEN_3644 : _GEN_3612; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3680 = _T_667 ? _GEN_3645 : _GEN_3613; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_3681 = _T_667 ? _GEN_3646 : _GEN_3614; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire  _GEN_3683 = _T_667 ? _GEN_2540 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_3691 = _T_637 ? _GEN_3647 : _GEN_2421; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3692 = _T_637 ? _GEN_2187 : _GEN_2422; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [6:0] _GEN_3693 = _T_637 ? _GEN_3649 : _GEN_2423; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3695 = _T_637 ? _GEN_3651 : _GEN_3584; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3696 = _T_637 ? _GEN_3652 : _GEN_3585; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3697 = _T_637 ? _GEN_3653 : _GEN_3586; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3698 = _T_637 ? _GEN_3654 : _GEN_3587; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3699 = _T_637 ? _GEN_3655 : _GEN_3588; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3700 = _T_637 ? _GEN_3656 : _GEN_3589; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3701 = _T_637 ? _GEN_3657 : _GEN_3590; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3702 = _T_637 ? _GEN_3658 : _GEN_3591; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3703 = _T_637 ? _GEN_3659 : _GEN_3592; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3704 = _T_637 ? _GEN_3660 : _GEN_3593; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3705 = _T_637 ? _GEN_3661 : _GEN_3594; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3706 = _T_637 ? _GEN_3662 : _GEN_3595; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3707 = _T_637 ? _GEN_3663 : _GEN_3596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3708 = _T_637 ? _GEN_3664 : _GEN_3597; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3709 = _T_637 ? _GEN_3665 : _GEN_3598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3710 = _T_637 ? _GEN_3666 : _GEN_3599; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3711 = _T_637 ? _GEN_3667 : _GEN_3600; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3712 = _T_637 ? _GEN_3668 : _GEN_3601; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3713 = _T_637 ? _GEN_3669 : _GEN_3602; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3714 = _T_637 ? _GEN_3670 : _GEN_3603; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3715 = _T_637 ? _GEN_3671 : _GEN_3604; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3716 = _T_637 ? _GEN_3672 : _GEN_3605; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3717 = _T_637 ? _GEN_3673 : _GEN_3606; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3718 = _T_637 ? _GEN_3674 : _GEN_3607; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3719 = _T_637 ? _GEN_3675 : _GEN_3608; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3720 = _T_637 ? _GEN_3676 : _GEN_3609; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3721 = _T_637 ? _GEN_3677 : _GEN_3610; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3722 = _T_637 ? _GEN_3678 : _GEN_3611; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3723 = _T_637 ? _GEN_3679 : _GEN_3612; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3724 = _T_637 ? _GEN_3680 : _GEN_3613; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3725 = _T_637 ? _GEN_3681 : _GEN_3614; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire  _GEN_3727 = _T_637 ? _GEN_3683 : _GEN_2540; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_3729 = 5'h1 == rd ? _next_reg_T_48 : _GEN_3695; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3730 = 5'h2 == rd ? _next_reg_T_48 : _GEN_3696; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3731 = 5'h3 == rd ? _next_reg_T_48 : _GEN_3697; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3732 = 5'h4 == rd ? _next_reg_T_48 : _GEN_3698; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3733 = 5'h5 == rd ? _next_reg_T_48 : _GEN_3699; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3734 = 5'h6 == rd ? _next_reg_T_48 : _GEN_3700; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3735 = 5'h7 == rd ? _next_reg_T_48 : _GEN_3701; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3736 = 5'h8 == rd ? _next_reg_T_48 : _GEN_3702; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3737 = 5'h9 == rd ? _next_reg_T_48 : _GEN_3703; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3738 = 5'ha == rd ? _next_reg_T_48 : _GEN_3704; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3739 = 5'hb == rd ? _next_reg_T_48 : _GEN_3705; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3740 = 5'hc == rd ? _next_reg_T_48 : _GEN_3706; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3741 = 5'hd == rd ? _next_reg_T_48 : _GEN_3707; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3742 = 5'he == rd ? _next_reg_T_48 : _GEN_3708; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3743 = 5'hf == rd ? _next_reg_T_48 : _GEN_3709; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3744 = 5'h10 == rd ? _next_reg_T_48 : _GEN_3710; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3745 = 5'h11 == rd ? _next_reg_T_48 : _GEN_3711; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3746 = 5'h12 == rd ? _next_reg_T_48 : _GEN_3712; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3747 = 5'h13 == rd ? _next_reg_T_48 : _GEN_3713; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3748 = 5'h14 == rd ? _next_reg_T_48 : _GEN_3714; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3749 = 5'h15 == rd ? _next_reg_T_48 : _GEN_3715; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3750 = 5'h16 == rd ? _next_reg_T_48 : _GEN_3716; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3751 = 5'h17 == rd ? _next_reg_T_48 : _GEN_3717; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3752 = 5'h18 == rd ? _next_reg_T_48 : _GEN_3718; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3753 = 5'h19 == rd ? _next_reg_T_48 : _GEN_3719; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3754 = 5'h1a == rd ? _next_reg_T_48 : _GEN_3720; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3755 = 5'h1b == rd ? _next_reg_T_48 : _GEN_3721; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3756 = 5'h1c == rd ? _next_reg_T_48 : _GEN_3722; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3757 = 5'h1d == rd ? _next_reg_T_48 : _GEN_3723; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3758 = 5'h1e == rd ? _next_reg_T_48 : _GEN_3724; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_3759 = 5'h1f == rd ? _next_reg_T_48 : _GEN_3725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire  _GEN_3760 = _T_669 | _GEN_3691; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [63:0] _GEN_3761 = _T_669 ? _T_663 : _T_663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55 423:23 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [6:0] _GEN_3762 = _T_669 ? 7'h40 : _GEN_3693; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [63:0] _GEN_3764 = _T_669 ? _GEN_3729 : _GEN_3695; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3765 = _T_669 ? _GEN_3730 : _GEN_3696; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3766 = _T_669 ? _GEN_3731 : _GEN_3697; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3767 = _T_669 ? _GEN_3732 : _GEN_3698; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3768 = _T_669 ? _GEN_3733 : _GEN_3699; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3769 = _T_669 ? _GEN_3734 : _GEN_3700; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3770 = _T_669 ? _GEN_3735 : _GEN_3701; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3771 = _T_669 ? _GEN_3736 : _GEN_3702; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3772 = _T_669 ? _GEN_3737 : _GEN_3703; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3773 = _T_669 ? _GEN_3738 : _GEN_3704; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3774 = _T_669 ? _GEN_3739 : _GEN_3705; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3775 = _T_669 ? _GEN_3740 : _GEN_3706; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3776 = _T_669 ? _GEN_3741 : _GEN_3707; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3777 = _T_669 ? _GEN_3742 : _GEN_3708; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3778 = _T_669 ? _GEN_3743 : _GEN_3709; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3779 = _T_669 ? _GEN_3744 : _GEN_3710; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3780 = _T_669 ? _GEN_3745 : _GEN_3711; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3781 = _T_669 ? _GEN_3746 : _GEN_3712; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3782 = _T_669 ? _GEN_3747 : _GEN_3713; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3783 = _T_669 ? _GEN_3748 : _GEN_3714; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3784 = _T_669 ? _GEN_3749 : _GEN_3715; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3785 = _T_669 ? _GEN_3750 : _GEN_3716; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3786 = _T_669 ? _GEN_3751 : _GEN_3717; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3787 = _T_669 ? _GEN_3752 : _GEN_3718; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3788 = _T_669 ? _GEN_3753 : _GEN_3719; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3789 = _T_669 ? _GEN_3754 : _GEN_3720; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3790 = _T_669 ? _GEN_3755 : _GEN_3721; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3791 = _T_669 ? _GEN_3756 : _GEN_3722; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3792 = _T_669 ? _GEN_3757 : _GEN_3723; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3793 = _T_669 ? _GEN_3758 : _GEN_3724; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_3794 = _T_669 ? _GEN_3759 : _GEN_3725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire  _GEN_3796 = _T_669 ? _GEN_3727 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_3804 = _T_657 ? _GEN_3760 : _GEN_3691; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3805 = _T_657 ? _GEN_3761 : _GEN_3692; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [6:0] _GEN_3806 = _T_657 ? _GEN_3762 : _GEN_3693; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3808 = _T_657 ? _GEN_3764 : _GEN_3695; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3809 = _T_657 ? _GEN_3765 : _GEN_3696; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3810 = _T_657 ? _GEN_3766 : _GEN_3697; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3811 = _T_657 ? _GEN_3767 : _GEN_3698; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3812 = _T_657 ? _GEN_3768 : _GEN_3699; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3813 = _T_657 ? _GEN_3769 : _GEN_3700; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3814 = _T_657 ? _GEN_3770 : _GEN_3701; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3815 = _T_657 ? _GEN_3771 : _GEN_3702; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3816 = _T_657 ? _GEN_3772 : _GEN_3703; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3817 = _T_657 ? _GEN_3773 : _GEN_3704; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3818 = _T_657 ? _GEN_3774 : _GEN_3705; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3819 = _T_657 ? _GEN_3775 : _GEN_3706; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3820 = _T_657 ? _GEN_3776 : _GEN_3707; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3821 = _T_657 ? _GEN_3777 : _GEN_3708; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3822 = _T_657 ? _GEN_3778 : _GEN_3709; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3823 = _T_657 ? _GEN_3779 : _GEN_3710; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3824 = _T_657 ? _GEN_3780 : _GEN_3711; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3825 = _T_657 ? _GEN_3781 : _GEN_3712; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3826 = _T_657 ? _GEN_3782 : _GEN_3713; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3827 = _T_657 ? _GEN_3783 : _GEN_3714; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3828 = _T_657 ? _GEN_3784 : _GEN_3715; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3829 = _T_657 ? _GEN_3785 : _GEN_3716; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3830 = _T_657 ? _GEN_3786 : _GEN_3717; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3831 = _T_657 ? _GEN_3787 : _GEN_3718; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3832 = _T_657 ? _GEN_3788 : _GEN_3719; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3833 = _T_657 ? _GEN_3789 : _GEN_3720; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3834 = _T_657 ? _GEN_3790 : _GEN_3721; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3835 = _T_657 ? _GEN_3791 : _GEN_3722; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3836 = _T_657 ? _GEN_3792 : _GEN_3723; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3837 = _T_657 ? _GEN_3793 : _GEN_3724; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_3838 = _T_657 ? _GEN_3794 : _GEN_3725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire  _GEN_3840 = _T_657 ? _GEN_3796 : _GEN_3727; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire  _GEN_3841 = _T_669 | _GEN_2508; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 82:26]
  wire [6:0] _GEN_3843 = _T_669 ? 7'h40 : _GEN_2510; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 84:26]
  wire [63:0] _GEN_3844 = _T_669 ? _GEN_840 : _GEN_2511; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:26]
  wire  _GEN_3846 = _T_669 ? _GEN_3840 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_3855 = _T_677 ? _GEN_3841 : _GEN_2508; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire [63:0] _GEN_3856 = _T_677 ? _GEN_3761 : _GEN_2509; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire [6:0] _GEN_3857 = _T_677 ? _GEN_3843 : _GEN_2510; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire [63:0] _GEN_3858 = _T_677 ? _GEN_3844 : _GEN_2511; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire  _GEN_3860 = _T_677 ? _GEN_3846 : _GEN_3840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire [63:0] _next_reg_T_176 = io_now_reg_2 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:52]
  wire [5:0] next_reg_rOff_7 = {_next_reg_T_176[2:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:48]
  wire [63:0] _next_reg_T_177 = io_mem_read_data >> next_reg_rOff_7; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:22]
  wire [63:0] _next_reg_T_178 = _next_reg_T_177 & 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire  next_reg_signBit_13 = _next_reg_T_178[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_181 = next_reg_signBit_13 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_182 = {_next_reg_T_181,_next_reg_T_178[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_3862 = 5'h1 == rd ? _next_reg_T_182 : _GEN_3808; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3863 = 5'h2 == rd ? _next_reg_T_182 : _GEN_3809; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3864 = 5'h3 == rd ? _next_reg_T_182 : _GEN_3810; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3865 = 5'h4 == rd ? _next_reg_T_182 : _GEN_3811; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3866 = 5'h5 == rd ? _next_reg_T_182 : _GEN_3812; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3867 = 5'h6 == rd ? _next_reg_T_182 : _GEN_3813; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3868 = 5'h7 == rd ? _next_reg_T_182 : _GEN_3814; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3869 = 5'h8 == rd ? _next_reg_T_182 : _GEN_3815; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3870 = 5'h9 == rd ? _next_reg_T_182 : _GEN_3816; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3871 = 5'ha == rd ? _next_reg_T_182 : _GEN_3817; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3872 = 5'hb == rd ? _next_reg_T_182 : _GEN_3818; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3873 = 5'hc == rd ? _next_reg_T_182 : _GEN_3819; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3874 = 5'hd == rd ? _next_reg_T_182 : _GEN_3820; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3875 = 5'he == rd ? _next_reg_T_182 : _GEN_3821; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3876 = 5'hf == rd ? _next_reg_T_182 : _GEN_3822; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3877 = 5'h10 == rd ? _next_reg_T_182 : _GEN_3823; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3878 = 5'h11 == rd ? _next_reg_T_182 : _GEN_3824; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3879 = 5'h12 == rd ? _next_reg_T_182 : _GEN_3825; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3880 = 5'h13 == rd ? _next_reg_T_182 : _GEN_3826; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3881 = 5'h14 == rd ? _next_reg_T_182 : _GEN_3827; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3882 = 5'h15 == rd ? _next_reg_T_182 : _GEN_3828; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3883 = 5'h16 == rd ? _next_reg_T_182 : _GEN_3829; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3884 = 5'h17 == rd ? _next_reg_T_182 : _GEN_3830; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3885 = 5'h18 == rd ? _next_reg_T_182 : _GEN_3831; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3886 = 5'h19 == rd ? _next_reg_T_182 : _GEN_3832; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3887 = 5'h1a == rd ? _next_reg_T_182 : _GEN_3833; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3888 = 5'h1b == rd ? _next_reg_T_182 : _GEN_3834; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3889 = 5'h1c == rd ? _next_reg_T_182 : _GEN_3835; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3890 = 5'h1d == rd ? _next_reg_T_182 : _GEN_3836; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3891 = 5'h1e == rd ? _next_reg_T_182 : _GEN_3837; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_3892 = 5'h1f == rd ? _next_reg_T_182 : _GEN_3838; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire  _GEN_3901 = _T_704 | _GEN_3804; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [63:0] _GEN_3902 = _T_704 ? _next_reg_T_176 : _GEN_3805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [6:0] _GEN_3903 = _T_704 ? 7'h20 : _GEN_3806; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [63:0] _GEN_3905 = _T_704 ? _GEN_3862 : _GEN_3808; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3906 = _T_704 ? _GEN_3863 : _GEN_3809; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3907 = _T_704 ? _GEN_3864 : _GEN_3810; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3908 = _T_704 ? _GEN_3865 : _GEN_3811; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3909 = _T_704 ? _GEN_3866 : _GEN_3812; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3910 = _T_704 ? _GEN_3867 : _GEN_3813; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3911 = _T_704 ? _GEN_3868 : _GEN_3814; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3912 = _T_704 ? _GEN_3869 : _GEN_3815; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3913 = _T_704 ? _GEN_3870 : _GEN_3816; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3914 = _T_704 ? _GEN_3871 : _GEN_3817; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3915 = _T_704 ? _GEN_3872 : _GEN_3818; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3916 = _T_704 ? _GEN_3873 : _GEN_3819; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3917 = _T_704 ? _GEN_3874 : _GEN_3820; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3918 = _T_704 ? _GEN_3875 : _GEN_3821; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3919 = _T_704 ? _GEN_3876 : _GEN_3822; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3920 = _T_704 ? _GEN_3877 : _GEN_3823; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3921 = _T_704 ? _GEN_3878 : _GEN_3824; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3922 = _T_704 ? _GEN_3879 : _GEN_3825; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3923 = _T_704 ? _GEN_3880 : _GEN_3826; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3924 = _T_704 ? _GEN_3881 : _GEN_3827; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3925 = _T_704 ? _GEN_3882 : _GEN_3828; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3926 = _T_704 ? _GEN_3883 : _GEN_3829; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3927 = _T_704 ? _GEN_3884 : _GEN_3830; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3928 = _T_704 ? _GEN_3885 : _GEN_3831; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3929 = _T_704 ? _GEN_3886 : _GEN_3832; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3930 = _T_704 ? _GEN_3887 : _GEN_3833; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3931 = _T_704 ? _GEN_3888 : _GEN_3834; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3932 = _T_704 ? _GEN_3889 : _GEN_3835; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3933 = _T_704 ? _GEN_3890 : _GEN_3836; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3934 = _T_704 ? _GEN_3891 : _GEN_3837; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_3935 = _T_704 ? _GEN_3892 : _GEN_3838; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire  _GEN_3942 = _T_711 | _GEN_3855; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 82:26]
  wire [63:0] _GEN_3943 = _T_711 ? _next_reg_T_176 : _GEN_3856; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 83:26]
  wire [6:0] _GEN_3944 = _T_711 ? 7'h20 : _GEN_3857; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 84:26]
  wire [63:0] _GEN_3945 = _T_711 ? {{32'd0}, _GEN_840[31:0]} : _GEN_3858; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:26]
  wire [2:0] _GEN_4013 = _T_720 ? inst[9:7] : 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 99:24]
  wire [2:0] _GEN_4120 = _T_729 ? inst[9:7] : _GEN_4013; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4198 = _T_770 ? inst[9:7] : _GEN_4120; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4242 = _T_779 ? inst[9:7] : _GEN_4198; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4711 = _T_875 ? inst[9:7] : _GEN_4242; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4815 = _T_889 ? inst[9:7] : _GEN_4711; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4919 = _T_897 ? inst[9:7] : _GEN_4815; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_5194 = _T_929 ? inst[9:7] : _GEN_4919; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_5329 = _T_937 ? inst[9:7] : _GEN_5194; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_5464 = _T_945 ? inst[9:7] : _GEN_5329; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_5599 = _T_953 ? inst[9:7] : _GEN_5464; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_5795 = _T_987 ? inst[9:7] : _GEN_5599; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_5902 = _T_996 ? inst[9:7] : _GEN_5795; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_6081 = _T_1018 ? inst[9:7] : _GEN_5902; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_6216 = _T_1026 ? inst[9:7] : _GEN_6081; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] rs1P = io_valid ? _GEN_6216 : 3'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 99:24]
  wire [2:0] _GEN_4015 = _T_720 ? inst[4:2] : 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 98:24]
  wire [2:0] _GEN_4201 = _T_770 ? rs1P : _GEN_4015; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:111 186:24]
  wire [2:0] _GEN_4245 = _T_779 ? rs1P : _GEN_4201; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:111 194:24]
  wire [2:0] _GEN_4538 = _T_846 ? inst[4:2] : _GEN_4245; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_4714 = _T_875 ? rs1P : _GEN_4538; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:111 235:24]
  wire [2:0] _GEN_4818 = _T_889 ? rs1P : _GEN_4714; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:111 240:24]
  wire [2:0] _GEN_4922 = _T_897 ? rs1P : _GEN_4818; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:111 245:24]
  wire [2:0] _GEN_5198 = _T_929 ? rs1P : _GEN_4922; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:111 253:23]
  wire [2:0] _GEN_5333 = _T_937 ? rs1P : _GEN_5198; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:111 254:23]
  wire [2:0] _GEN_5468 = _T_945 ? rs1P : _GEN_5333; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:111 255:23]
  wire [2:0] _GEN_5603 = _T_953 ? rs1P : _GEN_5468; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:111 256:23]
  wire [2:0] _GEN_5797 = _T_987 ? inst[4:2] : _GEN_5603; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_6085 = _T_1018 ? rs1P : _GEN_5797; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:111 297:24]
  wire [2:0] _GEN_6220 = _T_1026 ? rs1P : _GEN_6085; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:111 301:24]
  wire [2:0] rdP = io_valid ? _GEN_6220 : 3'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 98:24]
  wire [4:0] _T_727 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [4:0] _next_reg_T_183 = {2'h1,rs1P}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [63:0] _GEN_3947 = 5'h1 == _next_reg_T_183 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3948 = 5'h2 == _next_reg_T_183 ? io_now_reg_2 : _GEN_3947; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3949 = 5'h3 == _next_reg_T_183 ? io_now_reg_3 : _GEN_3948; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3950 = 5'h4 == _next_reg_T_183 ? io_now_reg_4 : _GEN_3949; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3951 = 5'h5 == _next_reg_T_183 ? io_now_reg_5 : _GEN_3950; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3952 = 5'h6 == _next_reg_T_183 ? io_now_reg_6 : _GEN_3951; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3953 = 5'h7 == _next_reg_T_183 ? io_now_reg_7 : _GEN_3952; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3954 = 5'h8 == _next_reg_T_183 ? io_now_reg_8 : _GEN_3953; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3955 = 5'h9 == _next_reg_T_183 ? io_now_reg_9 : _GEN_3954; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3956 = 5'ha == _next_reg_T_183 ? io_now_reg_10 : _GEN_3955; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3957 = 5'hb == _next_reg_T_183 ? io_now_reg_11 : _GEN_3956; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3958 = 5'hc == _next_reg_T_183 ? io_now_reg_12 : _GEN_3957; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3959 = 5'hd == _next_reg_T_183 ? io_now_reg_13 : _GEN_3958; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3960 = 5'he == _next_reg_T_183 ? io_now_reg_14 : _GEN_3959; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3961 = 5'hf == _next_reg_T_183 ? io_now_reg_15 : _GEN_3960; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3962 = 5'h10 == _next_reg_T_183 ? io_now_reg_16 : _GEN_3961; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3963 = 5'h11 == _next_reg_T_183 ? io_now_reg_17 : _GEN_3962; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3964 = 5'h12 == _next_reg_T_183 ? io_now_reg_18 : _GEN_3963; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3965 = 5'h13 == _next_reg_T_183 ? io_now_reg_19 : _GEN_3964; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3966 = 5'h14 == _next_reg_T_183 ? io_now_reg_20 : _GEN_3965; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3967 = 5'h15 == _next_reg_T_183 ? io_now_reg_21 : _GEN_3966; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3968 = 5'h16 == _next_reg_T_183 ? io_now_reg_22 : _GEN_3967; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3969 = 5'h17 == _next_reg_T_183 ? io_now_reg_23 : _GEN_3968; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3970 = 5'h18 == _next_reg_T_183 ? io_now_reg_24 : _GEN_3969; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3971 = 5'h19 == _next_reg_T_183 ? io_now_reg_25 : _GEN_3970; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3972 = 5'h1a == _next_reg_T_183 ? io_now_reg_26 : _GEN_3971; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3973 = 5'h1b == _next_reg_T_183 ? io_now_reg_27 : _GEN_3972; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3974 = 5'h1c == _next_reg_T_183 ? io_now_reg_28 : _GEN_3973; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3975 = 5'h1d == _next_reg_T_183 ? io_now_reg_29 : _GEN_3974; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3976 = 5'h1e == _next_reg_T_183 ? io_now_reg_30 : _GEN_3975; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_3977 = 5'h1f == _next_reg_T_183 ? io_now_reg_31 : _GEN_3976; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _next_reg_T_185 = _GEN_3977 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:68]
  wire [5:0] next_reg_rOff_8 = {_next_reg_T_185[2:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 50:48]
  wire [63:0] _next_reg_T_186 = io_mem_read_data >> next_reg_rOff_8; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:22]
  wire [63:0] _next_reg_T_187 = _next_reg_T_186 & 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 55:31]
  wire  next_reg_signBit_14 = _next_reg_T_187[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_190 = next_reg_signBit_14 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_191 = {_next_reg_T_190,_next_reg_T_187[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_3979 = 5'h1 == _T_727 ? _next_reg_T_191 : _GEN_3905; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3980 = 5'h2 == _T_727 ? _next_reg_T_191 : _GEN_3906; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3981 = 5'h3 == _T_727 ? _next_reg_T_191 : _GEN_3907; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3982 = 5'h4 == _T_727 ? _next_reg_T_191 : _GEN_3908; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3983 = 5'h5 == _T_727 ? _next_reg_T_191 : _GEN_3909; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3984 = 5'h6 == _T_727 ? _next_reg_T_191 : _GEN_3910; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3985 = 5'h7 == _T_727 ? _next_reg_T_191 : _GEN_3911; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3986 = 5'h8 == _T_727 ? _next_reg_T_191 : _GEN_3912; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3987 = 5'h9 == _T_727 ? _next_reg_T_191 : _GEN_3913; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3988 = 5'ha == _T_727 ? _next_reg_T_191 : _GEN_3914; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3989 = 5'hb == _T_727 ? _next_reg_T_191 : _GEN_3915; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3990 = 5'hc == _T_727 ? _next_reg_T_191 : _GEN_3916; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3991 = 5'hd == _T_727 ? _next_reg_T_191 : _GEN_3917; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3992 = 5'he == _T_727 ? _next_reg_T_191 : _GEN_3918; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3993 = 5'hf == _T_727 ? _next_reg_T_191 : _GEN_3919; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3994 = 5'h10 == _T_727 ? _next_reg_T_191 : _GEN_3920; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3995 = 5'h11 == _T_727 ? _next_reg_T_191 : _GEN_3921; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3996 = 5'h12 == _T_727 ? _next_reg_T_191 : _GEN_3922; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3997 = 5'h13 == _T_727 ? _next_reg_T_191 : _GEN_3923; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3998 = 5'h14 == _T_727 ? _next_reg_T_191 : _GEN_3924; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_3999 = 5'h15 == _T_727 ? _next_reg_T_191 : _GEN_3925; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_4000 = 5'h16 == _T_727 ? _next_reg_T_191 : _GEN_3926; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_4001 = 5'h17 == _T_727 ? _next_reg_T_191 : _GEN_3927; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_4002 = 5'h18 == _T_727 ? _next_reg_T_191 : _GEN_3928; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_4003 = 5'h19 == _T_727 ? _next_reg_T_191 : _GEN_3929; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_4004 = 5'h1a == _T_727 ? _next_reg_T_191 : _GEN_3930; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_4005 = 5'h1b == _T_727 ? _next_reg_T_191 : _GEN_3931; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_4006 = 5'h1c == _T_727 ? _next_reg_T_191 : _GEN_3932; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_4007 = 5'h1d == _T_727 ? _next_reg_T_191 : _GEN_3933; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_4008 = 5'h1e == _T_727 ? _next_reg_T_191 : _GEN_3934; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_4009 = 5'h1f == _T_727 ? _next_reg_T_191 : _GEN_3935; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire  _GEN_4018 = _T_720 | _GEN_3901; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [63:0] _GEN_4019 = _T_720 ? _next_reg_T_185 : _GEN_3902; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [6:0] _GEN_4020 = _T_720 ? 7'h20 : _GEN_3903; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [63:0] _GEN_4022 = _T_720 ? _GEN_3979 : _GEN_3905; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4023 = _T_720 ? _GEN_3980 : _GEN_3906; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4024 = _T_720 ? _GEN_3981 : _GEN_3907; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4025 = _T_720 ? _GEN_3982 : _GEN_3908; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4026 = _T_720 ? _GEN_3983 : _GEN_3909; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4027 = _T_720 ? _GEN_3984 : _GEN_3910; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4028 = _T_720 ? _GEN_3985 : _GEN_3911; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4029 = _T_720 ? _GEN_3986 : _GEN_3912; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4030 = _T_720 ? _GEN_3987 : _GEN_3913; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4031 = _T_720 ? _GEN_3988 : _GEN_3914; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4032 = _T_720 ? _GEN_3989 : _GEN_3915; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4033 = _T_720 ? _GEN_3990 : _GEN_3916; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4034 = _T_720 ? _GEN_3991 : _GEN_3917; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4035 = _T_720 ? _GEN_3992 : _GEN_3918; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4036 = _T_720 ? _GEN_3993 : _GEN_3919; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4037 = _T_720 ? _GEN_3994 : _GEN_3920; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4038 = _T_720 ? _GEN_3995 : _GEN_3921; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4039 = _T_720 ? _GEN_3996 : _GEN_3922; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4040 = _T_720 ? _GEN_3997 : _GEN_3923; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4041 = _T_720 ? _GEN_3998 : _GEN_3924; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4042 = _T_720 ? _GEN_3999 : _GEN_3925; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4043 = _T_720 ? _GEN_4000 : _GEN_3926; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4044 = _T_720 ? _GEN_4001 : _GEN_3927; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4045 = _T_720 ? _GEN_4002 : _GEN_3928; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4046 = _T_720 ? _GEN_4003 : _GEN_3929; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4047 = _T_720 ? _GEN_4004 : _GEN_3930; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4048 = _T_720 ? _GEN_4005 : _GEN_3931; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4049 = _T_720 ? _GEN_4006 : _GEN_3932; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4050 = _T_720 ? _GEN_4007 : _GEN_3933; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4051 = _T_720 ? _GEN_4008 : _GEN_3934; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_4052 = _T_720 ? _GEN_4009 : _GEN_3935; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [2:0] _GEN_4122 = _T_729 ? inst[4:2] : 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 100:24]
  wire [2:0] _GEN_5196 = _T_929 ? inst[4:2] : _GEN_4122; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_5331 = _T_937 ? inst[4:2] : _GEN_5196; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_5466 = _T_945 ? inst[4:2] : _GEN_5331; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_5601 = _T_953 ? inst[4:2] : _GEN_5466; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_5904 = _T_996 ? inst[4:2] : _GEN_5601; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_6083 = _T_1018 ? inst[4:2] : _GEN_5904; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_6218 = _T_1026 ? inst[4:2] : _GEN_6083; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] rs2P = io_valid ? _GEN_6218 : 3'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 100:24]
  wire [4:0] _T_739 = {2'h1,rs2P}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [63:0] _GEN_4086 = 5'h1 == _T_739 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4087 = 5'h2 == _T_739 ? io_now_reg_2 : _GEN_4086; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4088 = 5'h3 == _T_739 ? io_now_reg_3 : _GEN_4087; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4089 = 5'h4 == _T_739 ? io_now_reg_4 : _GEN_4088; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4090 = 5'h5 == _T_739 ? io_now_reg_5 : _GEN_4089; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4091 = 5'h6 == _T_739 ? io_now_reg_6 : _GEN_4090; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4092 = 5'h7 == _T_739 ? io_now_reg_7 : _GEN_4091; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4093 = 5'h8 == _T_739 ? io_now_reg_8 : _GEN_4092; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4094 = 5'h9 == _T_739 ? io_now_reg_9 : _GEN_4093; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4095 = 5'ha == _T_739 ? io_now_reg_10 : _GEN_4094; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4096 = 5'hb == _T_739 ? io_now_reg_11 : _GEN_4095; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4097 = 5'hc == _T_739 ? io_now_reg_12 : _GEN_4096; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4098 = 5'hd == _T_739 ? io_now_reg_13 : _GEN_4097; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4099 = 5'he == _T_739 ? io_now_reg_14 : _GEN_4098; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4100 = 5'hf == _T_739 ? io_now_reg_15 : _GEN_4099; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4101 = 5'h10 == _T_739 ? io_now_reg_16 : _GEN_4100; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4102 = 5'h11 == _T_739 ? io_now_reg_17 : _GEN_4101; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4103 = 5'h12 == _T_739 ? io_now_reg_18 : _GEN_4102; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4104 = 5'h13 == _T_739 ? io_now_reg_19 : _GEN_4103; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4105 = 5'h14 == _T_739 ? io_now_reg_20 : _GEN_4104; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4106 = 5'h15 == _T_739 ? io_now_reg_21 : _GEN_4105; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4107 = 5'h16 == _T_739 ? io_now_reg_22 : _GEN_4106; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4108 = 5'h17 == _T_739 ? io_now_reg_23 : _GEN_4107; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4109 = 5'h18 == _T_739 ? io_now_reg_24 : _GEN_4108; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4110 = 5'h19 == _T_739 ? io_now_reg_25 : _GEN_4109; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4111 = 5'h1a == _T_739 ? io_now_reg_26 : _GEN_4110; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4112 = 5'h1b == _T_739 ? io_now_reg_27 : _GEN_4111; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4113 = 5'h1c == _T_739 ? io_now_reg_28 : _GEN_4112; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4114 = 5'h1d == _T_739 ? io_now_reg_29 : _GEN_4113; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4115 = 5'h1e == _T_739 ? io_now_reg_30 : _GEN_4114; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire [63:0] _GEN_4116 = 5'h1f == _T_739 ? io_now_reg_31 : _GEN_4115; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:{26,26}]
  wire  _GEN_4125 = _T_729 | _GEN_3942; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 82:26]
  wire [63:0] _GEN_4126 = _T_729 ? _next_reg_T_185 : _GEN_3943; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 83:26]
  wire [6:0] _GEN_4127 = _T_729 ? 7'h20 : _GEN_3944; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 84:26]
  wire [63:0] _GEN_4128 = _T_729 ? _GEN_4116 : _GEN_3945; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:26]
  wire  _GEN_4134 = _T_741 | _GEN_1923; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 160:21 163:25]
  wire [63:0] _GEN_4135 = _T_741 ? _T_334 : _GEN_1924; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 160:21 164:25]
  wire [63:0] _next_reg_1_T_1 = io_now_pc + 64'h2; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 171:35]
  wire [63:0] _next_pc_T_23 = {_GEN_31[63:1],1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 177:21]
  wire  _GEN_4150 = _T_755 | _GEN_4134; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 175:25]
  wire [63:0] _GEN_4151 = _T_755 ? _next_pc_T_23 : _GEN_4135; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 177:15]
  wire  _GEN_4158 = _T_764 | _GEN_4150; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 181:25]
  wire [63:0] _GEN_4159 = _T_764 ? _next_pc_T_23 : _GEN_4151; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 183:21]
  wire [63:0] _GEN_4160 = _T_764 ? _next_reg_1_T_1 : _GEN_4022; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 184:21]
  wire  _GEN_4193 = _GEN_3977 == 64'h0 | _GEN_4158; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:42 190:27]
  wire [63:0] _GEN_4194 = _GEN_3977 == 64'h0 ? _T_334 : _GEN_4159; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:42 191:27]
  wire  _GEN_4203 = _T_770 ? _GEN_4193 : _GEN_4158; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24]
  wire [63:0] _GEN_4204 = _T_770 ? _GEN_4194 : _GEN_4159; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24]
  wire  _GEN_4237 = _GEN_3977 != 64'h0 | _GEN_4203; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:42 198:27]
  wire [63:0] _GEN_4238 = _GEN_3977 != 64'h0 ? _T_334 : _GEN_4204; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:42 199:27]
  wire  _GEN_4247 = _T_779 ? _GEN_4237 : _GEN_4203; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24]
  wire [63:0] _GEN_4248 = _T_779 ? _GEN_4238 : _GEN_4204; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24]
  wire [63:0] _GEN_4250 = 5'h1 == rd ? imm : _GEN_4160; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4251 = 5'h2 == rd ? imm : _GEN_4023; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4252 = 5'h3 == rd ? imm : _GEN_4024; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4253 = 5'h4 == rd ? imm : _GEN_4025; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4254 = 5'h5 == rd ? imm : _GEN_4026; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4255 = 5'h6 == rd ? imm : _GEN_4027; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4256 = 5'h7 == rd ? imm : _GEN_4028; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4257 = 5'h8 == rd ? imm : _GEN_4029; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4258 = 5'h9 == rd ? imm : _GEN_4030; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4259 = 5'ha == rd ? imm : _GEN_4031; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4260 = 5'hb == rd ? imm : _GEN_4032; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4261 = 5'hc == rd ? imm : _GEN_4033; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4262 = 5'hd == rd ? imm : _GEN_4034; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4263 = 5'he == rd ? imm : _GEN_4035; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4264 = 5'hf == rd ? imm : _GEN_4036; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4265 = 5'h10 == rd ? imm : _GEN_4037; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4266 = 5'h11 == rd ? imm : _GEN_4038; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4267 = 5'h12 == rd ? imm : _GEN_4039; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4268 = 5'h13 == rd ? imm : _GEN_4040; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4269 = 5'h14 == rd ? imm : _GEN_4041; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4270 = 5'h15 == rd ? imm : _GEN_4042; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4271 = 5'h16 == rd ? imm : _GEN_4043; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4272 = 5'h17 == rd ? imm : _GEN_4044; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4273 = 5'h18 == rd ? imm : _GEN_4045; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4274 = 5'h19 == rd ? imm : _GEN_4046; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4275 = 5'h1a == rd ? imm : _GEN_4047; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4276 = 5'h1b == rd ? imm : _GEN_4048; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4277 = 5'h1c == rd ? imm : _GEN_4049; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4278 = 5'h1d == rd ? imm : _GEN_4050; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4279 = 5'h1e == rd ? imm : _GEN_4051; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4280 = 5'h1f == rd ? imm : _GEN_4052; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_4290 = _T_791 ? _GEN_4250 : _GEN_4160; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4291 = _T_791 ? _GEN_4251 : _GEN_4023; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4292 = _T_791 ? _GEN_4252 : _GEN_4024; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4293 = _T_791 ? _GEN_4253 : _GEN_4025; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4294 = _T_791 ? _GEN_4254 : _GEN_4026; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4295 = _T_791 ? _GEN_4255 : _GEN_4027; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4296 = _T_791 ? _GEN_4256 : _GEN_4028; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4297 = _T_791 ? _GEN_4257 : _GEN_4029; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4298 = _T_791 ? _GEN_4258 : _GEN_4030; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4299 = _T_791 ? _GEN_4259 : _GEN_4031; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4300 = _T_791 ? _GEN_4260 : _GEN_4032; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4301 = _T_791 ? _GEN_4261 : _GEN_4033; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4302 = _T_791 ? _GEN_4262 : _GEN_4034; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4303 = _T_791 ? _GEN_4263 : _GEN_4035; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4304 = _T_791 ? _GEN_4264 : _GEN_4036; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4305 = _T_791 ? _GEN_4265 : _GEN_4037; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4306 = _T_791 ? _GEN_4266 : _GEN_4038; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4307 = _T_791 ? _GEN_4267 : _GEN_4039; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4308 = _T_791 ? _GEN_4268 : _GEN_4040; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4309 = _T_791 ? _GEN_4269 : _GEN_4041; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4310 = _T_791 ? _GEN_4270 : _GEN_4042; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4311 = _T_791 ? _GEN_4271 : _GEN_4043; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4312 = _T_791 ? _GEN_4272 : _GEN_4044; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4313 = _T_791 ? _GEN_4273 : _GEN_4045; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4314 = _T_791 ? _GEN_4274 : _GEN_4046; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4315 = _T_791 ? _GEN_4275 : _GEN_4047; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4316 = _T_791 ? _GEN_4276 : _GEN_4048; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4317 = _T_791 ? _GEN_4277 : _GEN_4049; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4318 = _T_791 ? _GEN_4278 : _GEN_4050; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4319 = _T_791 ? _GEN_4279 : _GEN_4051; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_4320 = _T_791 ? _GEN_4280 : _GEN_4052; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [17:0] _nzimm_C_LUI_T_7 = {inst[12],inst[6],inst[5],inst[4],inst[3],inst[2],12'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire  nzimm_C_LUI_signBit = _nzimm_C_LUI_T_7[17]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [45:0] _nzimm_C_LUI_T_9 = nzimm_C_LUI_signBit ? 46'h3fffffffffff : 46'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] nzimm_C_LUI = {_nzimm_C_LUI_T_9,inst[12],inst[6],inst[5],inst[4],inst[3],inst[2],12'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_4322 = 5'h1 == rd ? nzimm_C_LUI : _GEN_4290; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4323 = 5'h2 == rd ? nzimm_C_LUI : _GEN_4291; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4324 = 5'h3 == rd ? nzimm_C_LUI : _GEN_4292; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4325 = 5'h4 == rd ? nzimm_C_LUI : _GEN_4293; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4326 = 5'h5 == rd ? nzimm_C_LUI : _GEN_4294; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4327 = 5'h6 == rd ? nzimm_C_LUI : _GEN_4295; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4328 = 5'h7 == rd ? nzimm_C_LUI : _GEN_4296; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4329 = 5'h8 == rd ? nzimm_C_LUI : _GEN_4297; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4330 = 5'h9 == rd ? nzimm_C_LUI : _GEN_4298; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4331 = 5'ha == rd ? nzimm_C_LUI : _GEN_4299; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4332 = 5'hb == rd ? nzimm_C_LUI : _GEN_4300; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4333 = 5'hc == rd ? nzimm_C_LUI : _GEN_4301; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4334 = 5'hd == rd ? nzimm_C_LUI : _GEN_4302; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4335 = 5'he == rd ? nzimm_C_LUI : _GEN_4303; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4336 = 5'hf == rd ? nzimm_C_LUI : _GEN_4304; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4337 = 5'h10 == rd ? nzimm_C_LUI : _GEN_4305; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4338 = 5'h11 == rd ? nzimm_C_LUI : _GEN_4306; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4339 = 5'h12 == rd ? nzimm_C_LUI : _GEN_4307; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4340 = 5'h13 == rd ? nzimm_C_LUI : _GEN_4308; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4341 = 5'h14 == rd ? nzimm_C_LUI : _GEN_4309; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4342 = 5'h15 == rd ? nzimm_C_LUI : _GEN_4310; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4343 = 5'h16 == rd ? nzimm_C_LUI : _GEN_4311; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4344 = 5'h17 == rd ? nzimm_C_LUI : _GEN_4312; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4345 = 5'h18 == rd ? nzimm_C_LUI : _GEN_4313; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4346 = 5'h19 == rd ? nzimm_C_LUI : _GEN_4314; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4347 = 5'h1a == rd ? nzimm_C_LUI : _GEN_4315; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4348 = 5'h1b == rd ? nzimm_C_LUI : _GEN_4316; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4349 = 5'h1c == rd ? nzimm_C_LUI : _GEN_4317; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4350 = 5'h1d == rd ? nzimm_C_LUI : _GEN_4318; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4351 = 5'h1e == rd ? nzimm_C_LUI : _GEN_4319; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4352 = 5'h1f == rd ? nzimm_C_LUI : _GEN_4320; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_4361 = _T_809 ? _GEN_4322 : _GEN_4290; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4362 = _T_809 ? _GEN_4323 : _GEN_4291; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4363 = _T_809 ? _GEN_4324 : _GEN_4292; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4364 = _T_809 ? _GEN_4325 : _GEN_4293; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4365 = _T_809 ? _GEN_4326 : _GEN_4294; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4366 = _T_809 ? _GEN_4327 : _GEN_4295; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4367 = _T_809 ? _GEN_4328 : _GEN_4296; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4368 = _T_809 ? _GEN_4329 : _GEN_4297; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4369 = _T_809 ? _GEN_4330 : _GEN_4298; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4370 = _T_809 ? _GEN_4331 : _GEN_4299; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4371 = _T_809 ? _GEN_4332 : _GEN_4300; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4372 = _T_809 ? _GEN_4333 : _GEN_4301; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4373 = _T_809 ? _GEN_4334 : _GEN_4302; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4374 = _T_809 ? _GEN_4335 : _GEN_4303; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4375 = _T_809 ? _GEN_4336 : _GEN_4304; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4376 = _T_809 ? _GEN_4337 : _GEN_4305; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4377 = _T_809 ? _GEN_4338 : _GEN_4306; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4378 = _T_809 ? _GEN_4339 : _GEN_4307; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4379 = _T_809 ? _GEN_4340 : _GEN_4308; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4380 = _T_809 ? _GEN_4341 : _GEN_4309; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4381 = _T_809 ? _GEN_4342 : _GEN_4310; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4382 = _T_809 ? _GEN_4343 : _GEN_4311; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4383 = _T_809 ? _GEN_4344 : _GEN_4312; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4384 = _T_809 ? _GEN_4345 : _GEN_4313; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4385 = _T_809 ? _GEN_4346 : _GEN_4314; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4386 = _T_809 ? _GEN_4347 : _GEN_4315; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4387 = _T_809 ? _GEN_4348 : _GEN_4316; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4388 = _T_809 ? _GEN_4349 : _GEN_4317; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4389 = _T_809 ? _GEN_4350 : _GEN_4318; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4390 = _T_809 ? _GEN_4351 : _GEN_4319; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4391 = _T_809 ? _GEN_4352 : _GEN_4320; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_4393 = 5'h1 == rd ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4394 = 5'h2 == rd ? io_now_reg_2 : _GEN_4393; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4395 = 5'h3 == rd ? io_now_reg_3 : _GEN_4394; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4396 = 5'h4 == rd ? io_now_reg_4 : _GEN_4395; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4397 = 5'h5 == rd ? io_now_reg_5 : _GEN_4396; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4398 = 5'h6 == rd ? io_now_reg_6 : _GEN_4397; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4399 = 5'h7 == rd ? io_now_reg_7 : _GEN_4398; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4400 = 5'h8 == rd ? io_now_reg_8 : _GEN_4399; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4401 = 5'h9 == rd ? io_now_reg_9 : _GEN_4400; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4402 = 5'ha == rd ? io_now_reg_10 : _GEN_4401; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4403 = 5'hb == rd ? io_now_reg_11 : _GEN_4402; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4404 = 5'hc == rd ? io_now_reg_12 : _GEN_4403; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4405 = 5'hd == rd ? io_now_reg_13 : _GEN_4404; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4406 = 5'he == rd ? io_now_reg_14 : _GEN_4405; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4407 = 5'hf == rd ? io_now_reg_15 : _GEN_4406; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4408 = 5'h10 == rd ? io_now_reg_16 : _GEN_4407; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4409 = 5'h11 == rd ? io_now_reg_17 : _GEN_4408; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4410 = 5'h12 == rd ? io_now_reg_18 : _GEN_4409; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4411 = 5'h13 == rd ? io_now_reg_19 : _GEN_4410; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4412 = 5'h14 == rd ? io_now_reg_20 : _GEN_4411; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4413 = 5'h15 == rd ? io_now_reg_21 : _GEN_4412; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4414 = 5'h16 == rd ? io_now_reg_22 : _GEN_4413; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4415 = 5'h17 == rd ? io_now_reg_23 : _GEN_4414; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4416 = 5'h18 == rd ? io_now_reg_24 : _GEN_4415; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4417 = 5'h19 == rd ? io_now_reg_25 : _GEN_4416; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4418 = 5'h1a == rd ? io_now_reg_26 : _GEN_4417; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4419 = 5'h1b == rd ? io_now_reg_27 : _GEN_4418; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4420 = 5'h1c == rd ? io_now_reg_28 : _GEN_4419; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4421 = 5'h1d == rd ? io_now_reg_29 : _GEN_4420; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4422 = 5'h1e == rd ? io_now_reg_30 : _GEN_4421; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_4423 = 5'h1f == rd ? io_now_reg_31 : _GEN_4422; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _next_reg_T_193 = _GEN_4423 + _imm_T_309; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:35]
  wire [63:0] _GEN_4425 = 5'h1 == rd ? _next_reg_T_193 : _GEN_4361; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4426 = 5'h2 == rd ? _next_reg_T_193 : _GEN_4362; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4427 = 5'h3 == rd ? _next_reg_T_193 : _GEN_4363; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4428 = 5'h4 == rd ? _next_reg_T_193 : _GEN_4364; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4429 = 5'h5 == rd ? _next_reg_T_193 : _GEN_4365; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4430 = 5'h6 == rd ? _next_reg_T_193 : _GEN_4366; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4431 = 5'h7 == rd ? _next_reg_T_193 : _GEN_4367; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4432 = 5'h8 == rd ? _next_reg_T_193 : _GEN_4368; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4433 = 5'h9 == rd ? _next_reg_T_193 : _GEN_4369; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4434 = 5'ha == rd ? _next_reg_T_193 : _GEN_4370; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4435 = 5'hb == rd ? _next_reg_T_193 : _GEN_4371; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4436 = 5'hc == rd ? _next_reg_T_193 : _GEN_4372; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4437 = 5'hd == rd ? _next_reg_T_193 : _GEN_4373; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4438 = 5'he == rd ? _next_reg_T_193 : _GEN_4374; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4439 = 5'hf == rd ? _next_reg_T_193 : _GEN_4375; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4440 = 5'h10 == rd ? _next_reg_T_193 : _GEN_4376; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4441 = 5'h11 == rd ? _next_reg_T_193 : _GEN_4377; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4442 = 5'h12 == rd ? _next_reg_T_193 : _GEN_4378; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4443 = 5'h13 == rd ? _next_reg_T_193 : _GEN_4379; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4444 = 5'h14 == rd ? _next_reg_T_193 : _GEN_4380; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4445 = 5'h15 == rd ? _next_reg_T_193 : _GEN_4381; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4446 = 5'h16 == rd ? _next_reg_T_193 : _GEN_4382; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4447 = 5'h17 == rd ? _next_reg_T_193 : _GEN_4383; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4448 = 5'h18 == rd ? _next_reg_T_193 : _GEN_4384; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4449 = 5'h19 == rd ? _next_reg_T_193 : _GEN_4385; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4450 = 5'h1a == rd ? _next_reg_T_193 : _GEN_4386; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4451 = 5'h1b == rd ? _next_reg_T_193 : _GEN_4387; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4452 = 5'h1c == rd ? _next_reg_T_193 : _GEN_4388; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4453 = 5'h1d == rd ? _next_reg_T_193 : _GEN_4389; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4454 = 5'h1e == rd ? _next_reg_T_193 : _GEN_4390; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4455 = 5'h1f == rd ? _next_reg_T_193 : _GEN_4391; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_4464 = _T_824 ? _GEN_4425 : _GEN_4361; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4465 = _T_824 ? _GEN_4426 : _GEN_4362; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4466 = _T_824 ? _GEN_4427 : _GEN_4363; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4467 = _T_824 ? _GEN_4428 : _GEN_4364; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4468 = _T_824 ? _GEN_4429 : _GEN_4365; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4469 = _T_824 ? _GEN_4430 : _GEN_4366; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4470 = _T_824 ? _GEN_4431 : _GEN_4367; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4471 = _T_824 ? _GEN_4432 : _GEN_4368; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4472 = _T_824 ? _GEN_4433 : _GEN_4369; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4473 = _T_824 ? _GEN_4434 : _GEN_4370; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4474 = _T_824 ? _GEN_4435 : _GEN_4371; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4475 = _T_824 ? _GEN_4436 : _GEN_4372; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4476 = _T_824 ? _GEN_4437 : _GEN_4373; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4477 = _T_824 ? _GEN_4438 : _GEN_4374; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4478 = _T_824 ? _GEN_4439 : _GEN_4375; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4479 = _T_824 ? _GEN_4440 : _GEN_4376; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4480 = _T_824 ? _GEN_4441 : _GEN_4377; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4481 = _T_824 ? _GEN_4442 : _GEN_4378; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4482 = _T_824 ? _GEN_4443 : _GEN_4379; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4483 = _T_824 ? _GEN_4444 : _GEN_4380; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4484 = _T_824 ? _GEN_4445 : _GEN_4381; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4485 = _T_824 ? _GEN_4446 : _GEN_4382; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4486 = _T_824 ? _GEN_4447 : _GEN_4383; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4487 = _T_824 ? _GEN_4448 : _GEN_4384; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4488 = _T_824 ? _GEN_4449 : _GEN_4385; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4489 = _T_824 ? _GEN_4450 : _GEN_4386; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4490 = _T_824 ? _GEN_4451 : _GEN_4387; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4491 = _T_824 ? _GEN_4452 : _GEN_4388; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4492 = _T_824 ? _GEN_4453 : _GEN_4389; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4493 = _T_824 ? _GEN_4454 : _GEN_4390; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_4494 = _T_824 ? _GEN_4455 : _GEN_4391; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [9:0] _nzimm_C_ADDI16SP_T_7 = {inst[12],inst[4],inst[3],inst[5],inst[2],inst[6],4'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire  nzimm_C_ADDI16SP_signBit = _nzimm_C_ADDI16SP_T_7[9]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [53:0] _nzimm_C_ADDI16SP_T_9 = nzimm_C_ADDI16SP_signBit ? 54'h3fffffffffffff : 54'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] nzimm_C_ADDI16SP = {_nzimm_C_ADDI16SP_T_9,inst[12],inst[4],inst[3],inst[5],inst[2],inst[6],4'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _next_reg_2_T_1 = io_now_reg_2 + nzimm_C_ADDI16SP; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 223:37]
  wire [63:0] _GEN_4502 = _T_836 ? _next_reg_2_T_1 : _GEN_4465; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 220:28 223:21]
  wire [63:0] nzimm_C_ADDI4SPN = {54'h0,inst[10],inst[9],inst[8],inst[7],inst[12],inst[11],inst[5],inst[6],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [63:0] _next_reg_T_195 = io_now_reg_2 + nzimm_C_ADDI4SPN; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:44]
  wire [63:0] _GEN_4504 = 5'h1 == _T_727 ? _next_reg_T_195 : _GEN_4464; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4505 = 5'h2 == _T_727 ? _next_reg_T_195 : _GEN_4502; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4506 = 5'h3 == _T_727 ? _next_reg_T_195 : _GEN_4466; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4507 = 5'h4 == _T_727 ? _next_reg_T_195 : _GEN_4467; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4508 = 5'h5 == _T_727 ? _next_reg_T_195 : _GEN_4468; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4509 = 5'h6 == _T_727 ? _next_reg_T_195 : _GEN_4469; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4510 = 5'h7 == _T_727 ? _next_reg_T_195 : _GEN_4470; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4511 = 5'h8 == _T_727 ? _next_reg_T_195 : _GEN_4471; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4512 = 5'h9 == _T_727 ? _next_reg_T_195 : _GEN_4472; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4513 = 5'ha == _T_727 ? _next_reg_T_195 : _GEN_4473; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4514 = 5'hb == _T_727 ? _next_reg_T_195 : _GEN_4474; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4515 = 5'hc == _T_727 ? _next_reg_T_195 : _GEN_4475; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4516 = 5'hd == _T_727 ? _next_reg_T_195 : _GEN_4476; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4517 = 5'he == _T_727 ? _next_reg_T_195 : _GEN_4477; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4518 = 5'hf == _T_727 ? _next_reg_T_195 : _GEN_4478; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4519 = 5'h10 == _T_727 ? _next_reg_T_195 : _GEN_4479; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4520 = 5'h11 == _T_727 ? _next_reg_T_195 : _GEN_4480; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4521 = 5'h12 == _T_727 ? _next_reg_T_195 : _GEN_4481; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4522 = 5'h13 == _T_727 ? _next_reg_T_195 : _GEN_4482; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4523 = 5'h14 == _T_727 ? _next_reg_T_195 : _GEN_4483; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4524 = 5'h15 == _T_727 ? _next_reg_T_195 : _GEN_4484; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4525 = 5'h16 == _T_727 ? _next_reg_T_195 : _GEN_4485; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4526 = 5'h17 == _T_727 ? _next_reg_T_195 : _GEN_4486; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4527 = 5'h18 == _T_727 ? _next_reg_T_195 : _GEN_4487; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4528 = 5'h19 == _T_727 ? _next_reg_T_195 : _GEN_4488; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4529 = 5'h1a == _T_727 ? _next_reg_T_195 : _GEN_4489; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4530 = 5'h1b == _T_727 ? _next_reg_T_195 : _GEN_4490; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4531 = 5'h1c == _T_727 ? _next_reg_T_195 : _GEN_4491; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4532 = 5'h1d == _T_727 ? _next_reg_T_195 : _GEN_4492; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4533 = 5'h1e == _T_727 ? _next_reg_T_195 : _GEN_4493; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4534 = 5'h1f == _T_727 ? _next_reg_T_195 : _GEN_4494; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_4541 = _T_846 ? _GEN_4504 : _GEN_4464; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4542 = _T_846 ? _GEN_4505 : _GEN_4502; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4543 = _T_846 ? _GEN_4506 : _GEN_4466; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4544 = _T_846 ? _GEN_4507 : _GEN_4467; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4545 = _T_846 ? _GEN_4508 : _GEN_4468; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4546 = _T_846 ? _GEN_4509 : _GEN_4469; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4547 = _T_846 ? _GEN_4510 : _GEN_4470; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4548 = _T_846 ? _GEN_4511 : _GEN_4471; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4549 = _T_846 ? _GEN_4512 : _GEN_4472; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4550 = _T_846 ? _GEN_4513 : _GEN_4473; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4551 = _T_846 ? _GEN_4514 : _GEN_4474; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4552 = _T_846 ? _GEN_4515 : _GEN_4475; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4553 = _T_846 ? _GEN_4516 : _GEN_4476; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4554 = _T_846 ? _GEN_4517 : _GEN_4477; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4555 = _T_846 ? _GEN_4518 : _GEN_4478; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4556 = _T_846 ? _GEN_4519 : _GEN_4479; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4557 = _T_846 ? _GEN_4520 : _GEN_4480; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4558 = _T_846 ? _GEN_4521 : _GEN_4481; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4559 = _T_846 ? _GEN_4522 : _GEN_4482; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4560 = _T_846 ? _GEN_4523 : _GEN_4483; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4561 = _T_846 ? _GEN_4524 : _GEN_4484; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4562 = _T_846 ? _GEN_4525 : _GEN_4485; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4563 = _T_846 ? _GEN_4526 : _GEN_4486; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4564 = _T_846 ? _GEN_4527 : _GEN_4487; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4565 = _T_846 ? _GEN_4528 : _GEN_4488; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4566 = _T_846 ? _GEN_4529 : _GEN_4489; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4567 = _T_846 ? _GEN_4530 : _GEN_4490; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4568 = _T_846 ? _GEN_4531 : _GEN_4491; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4569 = _T_846 ? _GEN_4532 : _GEN_4492; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4570 = _T_846 ? _GEN_4533 : _GEN_4493; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_4571 = _T_846 ? _GEN_4534 : _GEN_4494; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [126:0] _GEN_138 = {{63'd0}, _GEN_4423}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:35]
  wire [126:0] _next_reg_T_197 = _GEN_138 << imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:35]
  wire [63:0] _GEN_4573 = 5'h1 == rd ? _next_reg_T_197[63:0] : _GEN_4541; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4574 = 5'h2 == rd ? _next_reg_T_197[63:0] : _GEN_4542; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4575 = 5'h3 == rd ? _next_reg_T_197[63:0] : _GEN_4543; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4576 = 5'h4 == rd ? _next_reg_T_197[63:0] : _GEN_4544; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4577 = 5'h5 == rd ? _next_reg_T_197[63:0] : _GEN_4545; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4578 = 5'h6 == rd ? _next_reg_T_197[63:0] : _GEN_4546; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4579 = 5'h7 == rd ? _next_reg_T_197[63:0] : _GEN_4547; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4580 = 5'h8 == rd ? _next_reg_T_197[63:0] : _GEN_4548; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4581 = 5'h9 == rd ? _next_reg_T_197[63:0] : _GEN_4549; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4582 = 5'ha == rd ? _next_reg_T_197[63:0] : _GEN_4550; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4583 = 5'hb == rd ? _next_reg_T_197[63:0] : _GEN_4551; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4584 = 5'hc == rd ? _next_reg_T_197[63:0] : _GEN_4552; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4585 = 5'hd == rd ? _next_reg_T_197[63:0] : _GEN_4553; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4586 = 5'he == rd ? _next_reg_T_197[63:0] : _GEN_4554; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4587 = 5'hf == rd ? _next_reg_T_197[63:0] : _GEN_4555; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4588 = 5'h10 == rd ? _next_reg_T_197[63:0] : _GEN_4556; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4589 = 5'h11 == rd ? _next_reg_T_197[63:0] : _GEN_4557; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4590 = 5'h12 == rd ? _next_reg_T_197[63:0] : _GEN_4558; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4591 = 5'h13 == rd ? _next_reg_T_197[63:0] : _GEN_4559; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4592 = 5'h14 == rd ? _next_reg_T_197[63:0] : _GEN_4560; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4593 = 5'h15 == rd ? _next_reg_T_197[63:0] : _GEN_4561; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4594 = 5'h16 == rd ? _next_reg_T_197[63:0] : _GEN_4562; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4595 = 5'h17 == rd ? _next_reg_T_197[63:0] : _GEN_4563; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4596 = 5'h18 == rd ? _next_reg_T_197[63:0] : _GEN_4564; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4597 = 5'h19 == rd ? _next_reg_T_197[63:0] : _GEN_4565; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4598 = 5'h1a == rd ? _next_reg_T_197[63:0] : _GEN_4566; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4599 = 5'h1b == rd ? _next_reg_T_197[63:0] : _GEN_4567; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4600 = 5'h1c == rd ? _next_reg_T_197[63:0] : _GEN_4568; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4601 = 5'h1d == rd ? _next_reg_T_197[63:0] : _GEN_4569; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4602 = 5'h1e == rd ? _next_reg_T_197[63:0] : _GEN_4570; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4603 = 5'h1f == rd ? _next_reg_T_197[63:0] : _GEN_4571; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_4613 = _T_862 ? _GEN_4573 : _GEN_4541; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4614 = _T_862 ? _GEN_4574 : _GEN_4542; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4615 = _T_862 ? _GEN_4575 : _GEN_4543; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4616 = _T_862 ? _GEN_4576 : _GEN_4544; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4617 = _T_862 ? _GEN_4577 : _GEN_4545; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4618 = _T_862 ? _GEN_4578 : _GEN_4546; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4619 = _T_862 ? _GEN_4579 : _GEN_4547; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4620 = _T_862 ? _GEN_4580 : _GEN_4548; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4621 = _T_862 ? _GEN_4581 : _GEN_4549; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4622 = _T_862 ? _GEN_4582 : _GEN_4550; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4623 = _T_862 ? _GEN_4583 : _GEN_4551; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4624 = _T_862 ? _GEN_4584 : _GEN_4552; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4625 = _T_862 ? _GEN_4585 : _GEN_4553; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4626 = _T_862 ? _GEN_4586 : _GEN_4554; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4627 = _T_862 ? _GEN_4587 : _GEN_4555; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4628 = _T_862 ? _GEN_4588 : _GEN_4556; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4629 = _T_862 ? _GEN_4589 : _GEN_4557; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4630 = _T_862 ? _GEN_4590 : _GEN_4558; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4631 = _T_862 ? _GEN_4591 : _GEN_4559; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4632 = _T_862 ? _GEN_4592 : _GEN_4560; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4633 = _T_862 ? _GEN_4593 : _GEN_4561; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4634 = _T_862 ? _GEN_4594 : _GEN_4562; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4635 = _T_862 ? _GEN_4595 : _GEN_4563; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4636 = _T_862 ? _GEN_4596 : _GEN_4564; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4637 = _T_862 ? _GEN_4597 : _GEN_4565; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4638 = _T_862 ? _GEN_4598 : _GEN_4566; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4639 = _T_862 ? _GEN_4599 : _GEN_4567; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4640 = _T_862 ? _GEN_4600 : _GEN_4568; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4641 = _T_862 ? _GEN_4601 : _GEN_4569; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4642 = _T_862 ? _GEN_4602 : _GEN_4570; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4643 = _T_862 ? _GEN_4603 : _GEN_4571; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_4645 = 5'h1 == _T_727 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4646 = 5'h2 == _T_727 ? io_now_reg_2 : _GEN_4645; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4647 = 5'h3 == _T_727 ? io_now_reg_3 : _GEN_4646; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4648 = 5'h4 == _T_727 ? io_now_reg_4 : _GEN_4647; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4649 = 5'h5 == _T_727 ? io_now_reg_5 : _GEN_4648; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4650 = 5'h6 == _T_727 ? io_now_reg_6 : _GEN_4649; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4651 = 5'h7 == _T_727 ? io_now_reg_7 : _GEN_4650; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4652 = 5'h8 == _T_727 ? io_now_reg_8 : _GEN_4651; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4653 = 5'h9 == _T_727 ? io_now_reg_9 : _GEN_4652; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4654 = 5'ha == _T_727 ? io_now_reg_10 : _GEN_4653; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4655 = 5'hb == _T_727 ? io_now_reg_11 : _GEN_4654; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4656 = 5'hc == _T_727 ? io_now_reg_12 : _GEN_4655; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4657 = 5'hd == _T_727 ? io_now_reg_13 : _GEN_4656; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4658 = 5'he == _T_727 ? io_now_reg_14 : _GEN_4657; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4659 = 5'hf == _T_727 ? io_now_reg_15 : _GEN_4658; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4660 = 5'h10 == _T_727 ? io_now_reg_16 : _GEN_4659; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4661 = 5'h11 == _T_727 ? io_now_reg_17 : _GEN_4660; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4662 = 5'h12 == _T_727 ? io_now_reg_18 : _GEN_4661; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4663 = 5'h13 == _T_727 ? io_now_reg_19 : _GEN_4662; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4664 = 5'h14 == _T_727 ? io_now_reg_20 : _GEN_4663; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4665 = 5'h15 == _T_727 ? io_now_reg_21 : _GEN_4664; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4666 = 5'h16 == _T_727 ? io_now_reg_22 : _GEN_4665; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4667 = 5'h17 == _T_727 ? io_now_reg_23 : _GEN_4666; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4668 = 5'h18 == _T_727 ? io_now_reg_24 : _GEN_4667; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4669 = 5'h19 == _T_727 ? io_now_reg_25 : _GEN_4668; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4670 = 5'h1a == _T_727 ? io_now_reg_26 : _GEN_4669; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4671 = 5'h1b == _T_727 ? io_now_reg_27 : _GEN_4670; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4672 = 5'h1c == _T_727 ? io_now_reg_28 : _GEN_4671; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4673 = 5'h1d == _T_727 ? io_now_reg_29 : _GEN_4672; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4674 = 5'h1e == _T_727 ? io_now_reg_30 : _GEN_4673; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_4675 = 5'h1f == _T_727 ? io_now_reg_31 : _GEN_4674; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _next_reg_T_200 = _GEN_4675 >> imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:51]
  wire [63:0] _GEN_4677 = 5'h1 == _T_727 ? _next_reg_T_200 : _GEN_4613; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4678 = 5'h2 == _T_727 ? _next_reg_T_200 : _GEN_4614; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4679 = 5'h3 == _T_727 ? _next_reg_T_200 : _GEN_4615; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4680 = 5'h4 == _T_727 ? _next_reg_T_200 : _GEN_4616; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4681 = 5'h5 == _T_727 ? _next_reg_T_200 : _GEN_4617; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4682 = 5'h6 == _T_727 ? _next_reg_T_200 : _GEN_4618; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4683 = 5'h7 == _T_727 ? _next_reg_T_200 : _GEN_4619; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4684 = 5'h8 == _T_727 ? _next_reg_T_200 : _GEN_4620; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4685 = 5'h9 == _T_727 ? _next_reg_T_200 : _GEN_4621; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4686 = 5'ha == _T_727 ? _next_reg_T_200 : _GEN_4622; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4687 = 5'hb == _T_727 ? _next_reg_T_200 : _GEN_4623; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4688 = 5'hc == _T_727 ? _next_reg_T_200 : _GEN_4624; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4689 = 5'hd == _T_727 ? _next_reg_T_200 : _GEN_4625; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4690 = 5'he == _T_727 ? _next_reg_T_200 : _GEN_4626; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4691 = 5'hf == _T_727 ? _next_reg_T_200 : _GEN_4627; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4692 = 5'h10 == _T_727 ? _next_reg_T_200 : _GEN_4628; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4693 = 5'h11 == _T_727 ? _next_reg_T_200 : _GEN_4629; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4694 = 5'h12 == _T_727 ? _next_reg_T_200 : _GEN_4630; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4695 = 5'h13 == _T_727 ? _next_reg_T_200 : _GEN_4631; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4696 = 5'h14 == _T_727 ? _next_reg_T_200 : _GEN_4632; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4697 = 5'h15 == _T_727 ? _next_reg_T_200 : _GEN_4633; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4698 = 5'h16 == _T_727 ? _next_reg_T_200 : _GEN_4634; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4699 = 5'h17 == _T_727 ? _next_reg_T_200 : _GEN_4635; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4700 = 5'h18 == _T_727 ? _next_reg_T_200 : _GEN_4636; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4701 = 5'h19 == _T_727 ? _next_reg_T_200 : _GEN_4637; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4702 = 5'h1a == _T_727 ? _next_reg_T_200 : _GEN_4638; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4703 = 5'h1b == _T_727 ? _next_reg_T_200 : _GEN_4639; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4704 = 5'h1c == _T_727 ? _next_reg_T_200 : _GEN_4640; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4705 = 5'h1d == _T_727 ? _next_reg_T_200 : _GEN_4641; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4706 = 5'h1e == _T_727 ? _next_reg_T_200 : _GEN_4642; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4707 = 5'h1f == _T_727 ? _next_reg_T_200 : _GEN_4643; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_4717 = _T_875 ? _GEN_4677 : _GEN_4613; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4718 = _T_875 ? _GEN_4678 : _GEN_4614; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4719 = _T_875 ? _GEN_4679 : _GEN_4615; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4720 = _T_875 ? _GEN_4680 : _GEN_4616; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4721 = _T_875 ? _GEN_4681 : _GEN_4617; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4722 = _T_875 ? _GEN_4682 : _GEN_4618; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4723 = _T_875 ? _GEN_4683 : _GEN_4619; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4724 = _T_875 ? _GEN_4684 : _GEN_4620; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4725 = _T_875 ? _GEN_4685 : _GEN_4621; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4726 = _T_875 ? _GEN_4686 : _GEN_4622; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4727 = _T_875 ? _GEN_4687 : _GEN_4623; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4728 = _T_875 ? _GEN_4688 : _GEN_4624; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4729 = _T_875 ? _GEN_4689 : _GEN_4625; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4730 = _T_875 ? _GEN_4690 : _GEN_4626; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4731 = _T_875 ? _GEN_4691 : _GEN_4627; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4732 = _T_875 ? _GEN_4692 : _GEN_4628; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4733 = _T_875 ? _GEN_4693 : _GEN_4629; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4734 = _T_875 ? _GEN_4694 : _GEN_4630; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4735 = _T_875 ? _GEN_4695 : _GEN_4631; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4736 = _T_875 ? _GEN_4696 : _GEN_4632; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4737 = _T_875 ? _GEN_4697 : _GEN_4633; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4738 = _T_875 ? _GEN_4698 : _GEN_4634; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4739 = _T_875 ? _GEN_4699 : _GEN_4635; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4740 = _T_875 ? _GEN_4700 : _GEN_4636; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4741 = _T_875 ? _GEN_4701 : _GEN_4637; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4742 = _T_875 ? _GEN_4702 : _GEN_4638; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4743 = _T_875 ? _GEN_4703 : _GEN_4639; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4744 = _T_875 ? _GEN_4704 : _GEN_4640; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4745 = _T_875 ? _GEN_4705 : _GEN_4641; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4746 = _T_875 ? _GEN_4706 : _GEN_4642; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_4747 = _T_875 ? _GEN_4707 : _GEN_4643; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _next_reg_T_202 = 5'h1f == _T_727 ? io_now_reg_31 : _GEN_4674; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:52]
  wire [63:0] _next_reg_T_205 = $signed(_next_reg_T_202) >>> imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:73]
  wire [63:0] _GEN_4781 = 5'h1 == _T_727 ? _next_reg_T_205 : _GEN_4717; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4782 = 5'h2 == _T_727 ? _next_reg_T_205 : _GEN_4718; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4783 = 5'h3 == _T_727 ? _next_reg_T_205 : _GEN_4719; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4784 = 5'h4 == _T_727 ? _next_reg_T_205 : _GEN_4720; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4785 = 5'h5 == _T_727 ? _next_reg_T_205 : _GEN_4721; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4786 = 5'h6 == _T_727 ? _next_reg_T_205 : _GEN_4722; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4787 = 5'h7 == _T_727 ? _next_reg_T_205 : _GEN_4723; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4788 = 5'h8 == _T_727 ? _next_reg_T_205 : _GEN_4724; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4789 = 5'h9 == _T_727 ? _next_reg_T_205 : _GEN_4725; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4790 = 5'ha == _T_727 ? _next_reg_T_205 : _GEN_4726; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4791 = 5'hb == _T_727 ? _next_reg_T_205 : _GEN_4727; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4792 = 5'hc == _T_727 ? _next_reg_T_205 : _GEN_4728; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4793 = 5'hd == _T_727 ? _next_reg_T_205 : _GEN_4729; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4794 = 5'he == _T_727 ? _next_reg_T_205 : _GEN_4730; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4795 = 5'hf == _T_727 ? _next_reg_T_205 : _GEN_4731; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4796 = 5'h10 == _T_727 ? _next_reg_T_205 : _GEN_4732; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4797 = 5'h11 == _T_727 ? _next_reg_T_205 : _GEN_4733; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4798 = 5'h12 == _T_727 ? _next_reg_T_205 : _GEN_4734; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4799 = 5'h13 == _T_727 ? _next_reg_T_205 : _GEN_4735; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4800 = 5'h14 == _T_727 ? _next_reg_T_205 : _GEN_4736; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4801 = 5'h15 == _T_727 ? _next_reg_T_205 : _GEN_4737; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4802 = 5'h16 == _T_727 ? _next_reg_T_205 : _GEN_4738; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4803 = 5'h17 == _T_727 ? _next_reg_T_205 : _GEN_4739; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4804 = 5'h18 == _T_727 ? _next_reg_T_205 : _GEN_4740; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4805 = 5'h19 == _T_727 ? _next_reg_T_205 : _GEN_4741; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4806 = 5'h1a == _T_727 ? _next_reg_T_205 : _GEN_4742; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4807 = 5'h1b == _T_727 ? _next_reg_T_205 : _GEN_4743; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4808 = 5'h1c == _T_727 ? _next_reg_T_205 : _GEN_4744; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4809 = 5'h1d == _T_727 ? _next_reg_T_205 : _GEN_4745; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4810 = 5'h1e == _T_727 ? _next_reg_T_205 : _GEN_4746; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4811 = 5'h1f == _T_727 ? _next_reg_T_205 : _GEN_4747; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_4821 = _T_889 ? _GEN_4781 : _GEN_4717; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4822 = _T_889 ? _GEN_4782 : _GEN_4718; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4823 = _T_889 ? _GEN_4783 : _GEN_4719; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4824 = _T_889 ? _GEN_4784 : _GEN_4720; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4825 = _T_889 ? _GEN_4785 : _GEN_4721; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4826 = _T_889 ? _GEN_4786 : _GEN_4722; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4827 = _T_889 ? _GEN_4787 : _GEN_4723; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4828 = _T_889 ? _GEN_4788 : _GEN_4724; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4829 = _T_889 ? _GEN_4789 : _GEN_4725; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4830 = _T_889 ? _GEN_4790 : _GEN_4726; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4831 = _T_889 ? _GEN_4791 : _GEN_4727; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4832 = _T_889 ? _GEN_4792 : _GEN_4728; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4833 = _T_889 ? _GEN_4793 : _GEN_4729; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4834 = _T_889 ? _GEN_4794 : _GEN_4730; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4835 = _T_889 ? _GEN_4795 : _GEN_4731; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4836 = _T_889 ? _GEN_4796 : _GEN_4732; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4837 = _T_889 ? _GEN_4797 : _GEN_4733; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4838 = _T_889 ? _GEN_4798 : _GEN_4734; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4839 = _T_889 ? _GEN_4799 : _GEN_4735; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4840 = _T_889 ? _GEN_4800 : _GEN_4736; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4841 = _T_889 ? _GEN_4801 : _GEN_4737; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4842 = _T_889 ? _GEN_4802 : _GEN_4738; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4843 = _T_889 ? _GEN_4803 : _GEN_4739; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4844 = _T_889 ? _GEN_4804 : _GEN_4740; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4845 = _T_889 ? _GEN_4805 : _GEN_4741; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4846 = _T_889 ? _GEN_4806 : _GEN_4742; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4847 = _T_889 ? _GEN_4807 : _GEN_4743; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4848 = _T_889 ? _GEN_4808 : _GEN_4744; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4849 = _T_889 ? _GEN_4809 : _GEN_4745; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4850 = _T_889 ? _GEN_4810 : _GEN_4746; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_4851 = _T_889 ? _GEN_4811 : _GEN_4747; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _next_reg_T_207 = _GEN_4675 & imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:51]
  wire [63:0] _GEN_4885 = 5'h1 == _T_727 ? _next_reg_T_207 : _GEN_4821; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4886 = 5'h2 == _T_727 ? _next_reg_T_207 : _GEN_4822; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4887 = 5'h3 == _T_727 ? _next_reg_T_207 : _GEN_4823; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4888 = 5'h4 == _T_727 ? _next_reg_T_207 : _GEN_4824; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4889 = 5'h5 == _T_727 ? _next_reg_T_207 : _GEN_4825; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4890 = 5'h6 == _T_727 ? _next_reg_T_207 : _GEN_4826; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4891 = 5'h7 == _T_727 ? _next_reg_T_207 : _GEN_4827; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4892 = 5'h8 == _T_727 ? _next_reg_T_207 : _GEN_4828; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4893 = 5'h9 == _T_727 ? _next_reg_T_207 : _GEN_4829; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4894 = 5'ha == _T_727 ? _next_reg_T_207 : _GEN_4830; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4895 = 5'hb == _T_727 ? _next_reg_T_207 : _GEN_4831; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4896 = 5'hc == _T_727 ? _next_reg_T_207 : _GEN_4832; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4897 = 5'hd == _T_727 ? _next_reg_T_207 : _GEN_4833; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4898 = 5'he == _T_727 ? _next_reg_T_207 : _GEN_4834; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4899 = 5'hf == _T_727 ? _next_reg_T_207 : _GEN_4835; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4900 = 5'h10 == _T_727 ? _next_reg_T_207 : _GEN_4836; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4901 = 5'h11 == _T_727 ? _next_reg_T_207 : _GEN_4837; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4902 = 5'h12 == _T_727 ? _next_reg_T_207 : _GEN_4838; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4903 = 5'h13 == _T_727 ? _next_reg_T_207 : _GEN_4839; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4904 = 5'h14 == _T_727 ? _next_reg_T_207 : _GEN_4840; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4905 = 5'h15 == _T_727 ? _next_reg_T_207 : _GEN_4841; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4906 = 5'h16 == _T_727 ? _next_reg_T_207 : _GEN_4842; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4907 = 5'h17 == _T_727 ? _next_reg_T_207 : _GEN_4843; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4908 = 5'h18 == _T_727 ? _next_reg_T_207 : _GEN_4844; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4909 = 5'h19 == _T_727 ? _next_reg_T_207 : _GEN_4845; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4910 = 5'h1a == _T_727 ? _next_reg_T_207 : _GEN_4846; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4911 = 5'h1b == _T_727 ? _next_reg_T_207 : _GEN_4847; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4912 = 5'h1c == _T_727 ? _next_reg_T_207 : _GEN_4848; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4913 = 5'h1d == _T_727 ? _next_reg_T_207 : _GEN_4849; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4914 = 5'h1e == _T_727 ? _next_reg_T_207 : _GEN_4850; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4915 = 5'h1f == _T_727 ? _next_reg_T_207 : _GEN_4851; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_4925 = _T_897 ? _GEN_4885 : _GEN_4821; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4926 = _T_897 ? _GEN_4886 : _GEN_4822; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4927 = _T_897 ? _GEN_4887 : _GEN_4823; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4928 = _T_897 ? _GEN_4888 : _GEN_4824; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4929 = _T_897 ? _GEN_4889 : _GEN_4825; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4930 = _T_897 ? _GEN_4890 : _GEN_4826; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4931 = _T_897 ? _GEN_4891 : _GEN_4827; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4932 = _T_897 ? _GEN_4892 : _GEN_4828; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4933 = _T_897 ? _GEN_4893 : _GEN_4829; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4934 = _T_897 ? _GEN_4894 : _GEN_4830; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4935 = _T_897 ? _GEN_4895 : _GEN_4831; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4936 = _T_897 ? _GEN_4896 : _GEN_4832; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4937 = _T_897 ? _GEN_4897 : _GEN_4833; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4938 = _T_897 ? _GEN_4898 : _GEN_4834; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4939 = _T_897 ? _GEN_4899 : _GEN_4835; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4940 = _T_897 ? _GEN_4900 : _GEN_4836; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4941 = _T_897 ? _GEN_4901 : _GEN_4837; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4942 = _T_897 ? _GEN_4902 : _GEN_4838; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4943 = _T_897 ? _GEN_4903 : _GEN_4839; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4944 = _T_897 ? _GEN_4904 : _GEN_4840; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4945 = _T_897 ? _GEN_4905 : _GEN_4841; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4946 = _T_897 ? _GEN_4906 : _GEN_4842; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4947 = _T_897 ? _GEN_4907 : _GEN_4843; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4948 = _T_897 ? _GEN_4908 : _GEN_4844; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4949 = _T_897 ? _GEN_4909 : _GEN_4845; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4950 = _T_897 ? _GEN_4910 : _GEN_4846; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4951 = _T_897 ? _GEN_4911 : _GEN_4847; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4952 = _T_897 ? _GEN_4912 : _GEN_4848; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4953 = _T_897 ? _GEN_4913 : _GEN_4849; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4954 = _T_897 ? _GEN_4914 : _GEN_4850; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_4955 = _T_897 ? _GEN_4915 : _GEN_4851; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _next_reg_T_209 = io_now_reg_0 + _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:64]
  wire [63:0] _GEN_4957 = 5'h1 == rd ? _next_reg_T_209 : _GEN_4925; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4958 = 5'h2 == rd ? _next_reg_T_209 : _GEN_4926; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4959 = 5'h3 == rd ? _next_reg_T_209 : _GEN_4927; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4960 = 5'h4 == rd ? _next_reg_T_209 : _GEN_4928; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4961 = 5'h5 == rd ? _next_reg_T_209 : _GEN_4929; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4962 = 5'h6 == rd ? _next_reg_T_209 : _GEN_4930; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4963 = 5'h7 == rd ? _next_reg_T_209 : _GEN_4931; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4964 = 5'h8 == rd ? _next_reg_T_209 : _GEN_4932; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4965 = 5'h9 == rd ? _next_reg_T_209 : _GEN_4933; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4966 = 5'ha == rd ? _next_reg_T_209 : _GEN_4934; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4967 = 5'hb == rd ? _next_reg_T_209 : _GEN_4935; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4968 = 5'hc == rd ? _next_reg_T_209 : _GEN_4936; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4969 = 5'hd == rd ? _next_reg_T_209 : _GEN_4937; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4970 = 5'he == rd ? _next_reg_T_209 : _GEN_4938; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4971 = 5'hf == rd ? _next_reg_T_209 : _GEN_4939; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4972 = 5'h10 == rd ? _next_reg_T_209 : _GEN_4940; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4973 = 5'h11 == rd ? _next_reg_T_209 : _GEN_4941; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4974 = 5'h12 == rd ? _next_reg_T_209 : _GEN_4942; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4975 = 5'h13 == rd ? _next_reg_T_209 : _GEN_4943; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4976 = 5'h14 == rd ? _next_reg_T_209 : _GEN_4944; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4977 = 5'h15 == rd ? _next_reg_T_209 : _GEN_4945; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4978 = 5'h16 == rd ? _next_reg_T_209 : _GEN_4946; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4979 = 5'h17 == rd ? _next_reg_T_209 : _GEN_4947; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4980 = 5'h18 == rd ? _next_reg_T_209 : _GEN_4948; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4981 = 5'h19 == rd ? _next_reg_T_209 : _GEN_4949; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4982 = 5'h1a == rd ? _next_reg_T_209 : _GEN_4950; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4983 = 5'h1b == rd ? _next_reg_T_209 : _GEN_4951; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4984 = 5'h1c == rd ? _next_reg_T_209 : _GEN_4952; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4985 = 5'h1d == rd ? _next_reg_T_209 : _GEN_4953; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4986 = 5'h1e == rd ? _next_reg_T_209 : _GEN_4954; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4987 = 5'h1f == rd ? _next_reg_T_209 : _GEN_4955; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_4995 = _T_911 ? _GEN_4957 : _GEN_4925; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_4996 = _T_911 ? _GEN_4958 : _GEN_4926; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_4997 = _T_911 ? _GEN_4959 : _GEN_4927; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_4998 = _T_911 ? _GEN_4960 : _GEN_4928; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_4999 = _T_911 ? _GEN_4961 : _GEN_4929; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5000 = _T_911 ? _GEN_4962 : _GEN_4930; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5001 = _T_911 ? _GEN_4963 : _GEN_4931; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5002 = _T_911 ? _GEN_4964 : _GEN_4932; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5003 = _T_911 ? _GEN_4965 : _GEN_4933; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5004 = _T_911 ? _GEN_4966 : _GEN_4934; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5005 = _T_911 ? _GEN_4967 : _GEN_4935; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5006 = _T_911 ? _GEN_4968 : _GEN_4936; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5007 = _T_911 ? _GEN_4969 : _GEN_4937; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5008 = _T_911 ? _GEN_4970 : _GEN_4938; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5009 = _T_911 ? _GEN_4971 : _GEN_4939; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5010 = _T_911 ? _GEN_4972 : _GEN_4940; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5011 = _T_911 ? _GEN_4973 : _GEN_4941; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5012 = _T_911 ? _GEN_4974 : _GEN_4942; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5013 = _T_911 ? _GEN_4975 : _GEN_4943; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5014 = _T_911 ? _GEN_4976 : _GEN_4944; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5015 = _T_911 ? _GEN_4977 : _GEN_4945; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5016 = _T_911 ? _GEN_4978 : _GEN_4946; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5017 = _T_911 ? _GEN_4979 : _GEN_4947; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5018 = _T_911 ? _GEN_4980 : _GEN_4948; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5019 = _T_911 ? _GEN_4981 : _GEN_4949; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5020 = _T_911 ? _GEN_4982 : _GEN_4950; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5021 = _T_911 ? _GEN_4983 : _GEN_4951; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5022 = _T_911 ? _GEN_4984 : _GEN_4952; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5023 = _T_911 ? _GEN_4985 : _GEN_4953; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5024 = _T_911 ? _GEN_4986 : _GEN_4954; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_5025 = _T_911 ? _GEN_4987 : _GEN_4955; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _next_reg_T_211 = _GEN_4423 + _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:63]
  wire [63:0] _GEN_5027 = 5'h1 == rd ? _next_reg_T_211 : _GEN_4995; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5028 = 5'h2 == rd ? _next_reg_T_211 : _GEN_4996; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5029 = 5'h3 == rd ? _next_reg_T_211 : _GEN_4997; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5030 = 5'h4 == rd ? _next_reg_T_211 : _GEN_4998; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5031 = 5'h5 == rd ? _next_reg_T_211 : _GEN_4999; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5032 = 5'h6 == rd ? _next_reg_T_211 : _GEN_5000; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5033 = 5'h7 == rd ? _next_reg_T_211 : _GEN_5001; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5034 = 5'h8 == rd ? _next_reg_T_211 : _GEN_5002; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5035 = 5'h9 == rd ? _next_reg_T_211 : _GEN_5003; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5036 = 5'ha == rd ? _next_reg_T_211 : _GEN_5004; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5037 = 5'hb == rd ? _next_reg_T_211 : _GEN_5005; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5038 = 5'hc == rd ? _next_reg_T_211 : _GEN_5006; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5039 = 5'hd == rd ? _next_reg_T_211 : _GEN_5007; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5040 = 5'he == rd ? _next_reg_T_211 : _GEN_5008; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5041 = 5'hf == rd ? _next_reg_T_211 : _GEN_5009; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5042 = 5'h10 == rd ? _next_reg_T_211 : _GEN_5010; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5043 = 5'h11 == rd ? _next_reg_T_211 : _GEN_5011; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5044 = 5'h12 == rd ? _next_reg_T_211 : _GEN_5012; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5045 = 5'h13 == rd ? _next_reg_T_211 : _GEN_5013; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5046 = 5'h14 == rd ? _next_reg_T_211 : _GEN_5014; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5047 = 5'h15 == rd ? _next_reg_T_211 : _GEN_5015; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5048 = 5'h16 == rd ? _next_reg_T_211 : _GEN_5016; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5049 = 5'h17 == rd ? _next_reg_T_211 : _GEN_5017; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5050 = 5'h18 == rd ? _next_reg_T_211 : _GEN_5018; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5051 = 5'h19 == rd ? _next_reg_T_211 : _GEN_5019; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5052 = 5'h1a == rd ? _next_reg_T_211 : _GEN_5020; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5053 = 5'h1b == rd ? _next_reg_T_211 : _GEN_5021; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5054 = 5'h1c == rd ? _next_reg_T_211 : _GEN_5022; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5055 = 5'h1d == rd ? _next_reg_T_211 : _GEN_5023; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5056 = 5'h1e == rd ? _next_reg_T_211 : _GEN_5024; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5057 = 5'h1f == rd ? _next_reg_T_211 : _GEN_5025; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_5065 = _T_923 ? _GEN_5027 : _GEN_4995; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5066 = _T_923 ? _GEN_5028 : _GEN_4996; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5067 = _T_923 ? _GEN_5029 : _GEN_4997; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5068 = _T_923 ? _GEN_5030 : _GEN_4998; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5069 = _T_923 ? _GEN_5031 : _GEN_4999; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5070 = _T_923 ? _GEN_5032 : _GEN_5000; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5071 = _T_923 ? _GEN_5033 : _GEN_5001; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5072 = _T_923 ? _GEN_5034 : _GEN_5002; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5073 = _T_923 ? _GEN_5035 : _GEN_5003; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5074 = _T_923 ? _GEN_5036 : _GEN_5004; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5075 = _T_923 ? _GEN_5037 : _GEN_5005; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5076 = _T_923 ? _GEN_5038 : _GEN_5006; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5077 = _T_923 ? _GEN_5039 : _GEN_5007; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5078 = _T_923 ? _GEN_5040 : _GEN_5008; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5079 = _T_923 ? _GEN_5041 : _GEN_5009; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5080 = _T_923 ? _GEN_5042 : _GEN_5010; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5081 = _T_923 ? _GEN_5043 : _GEN_5011; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5082 = _T_923 ? _GEN_5044 : _GEN_5012; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5083 = _T_923 ? _GEN_5045 : _GEN_5013; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5084 = _T_923 ? _GEN_5046 : _GEN_5014; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5085 = _T_923 ? _GEN_5047 : _GEN_5015; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5086 = _T_923 ? _GEN_5048 : _GEN_5016; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5087 = _T_923 ? _GEN_5049 : _GEN_5017; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5088 = _T_923 ? _GEN_5050 : _GEN_5018; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5089 = _T_923 ? _GEN_5051 : _GEN_5019; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5090 = _T_923 ? _GEN_5052 : _GEN_5020; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5091 = _T_923 ? _GEN_5053 : _GEN_5021; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5092 = _T_923 ? _GEN_5054 : _GEN_5022; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5093 = _T_923 ? _GEN_5055 : _GEN_5023; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5094 = _T_923 ? _GEN_5056 : _GEN_5024; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_5095 = _T_923 ? _GEN_5057 : _GEN_5025; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _next_reg_T_214 = _GEN_4675 & _GEN_4116; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:79]
  wire [63:0] _GEN_5161 = 5'h1 == _T_727 ? _next_reg_T_214 : _GEN_5065; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5162 = 5'h2 == _T_727 ? _next_reg_T_214 : _GEN_5066; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5163 = 5'h3 == _T_727 ? _next_reg_T_214 : _GEN_5067; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5164 = 5'h4 == _T_727 ? _next_reg_T_214 : _GEN_5068; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5165 = 5'h5 == _T_727 ? _next_reg_T_214 : _GEN_5069; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5166 = 5'h6 == _T_727 ? _next_reg_T_214 : _GEN_5070; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5167 = 5'h7 == _T_727 ? _next_reg_T_214 : _GEN_5071; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5168 = 5'h8 == _T_727 ? _next_reg_T_214 : _GEN_5072; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5169 = 5'h9 == _T_727 ? _next_reg_T_214 : _GEN_5073; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5170 = 5'ha == _T_727 ? _next_reg_T_214 : _GEN_5074; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5171 = 5'hb == _T_727 ? _next_reg_T_214 : _GEN_5075; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5172 = 5'hc == _T_727 ? _next_reg_T_214 : _GEN_5076; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5173 = 5'hd == _T_727 ? _next_reg_T_214 : _GEN_5077; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5174 = 5'he == _T_727 ? _next_reg_T_214 : _GEN_5078; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5175 = 5'hf == _T_727 ? _next_reg_T_214 : _GEN_5079; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5176 = 5'h10 == _T_727 ? _next_reg_T_214 : _GEN_5080; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5177 = 5'h11 == _T_727 ? _next_reg_T_214 : _GEN_5081; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5178 = 5'h12 == _T_727 ? _next_reg_T_214 : _GEN_5082; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5179 = 5'h13 == _T_727 ? _next_reg_T_214 : _GEN_5083; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5180 = 5'h14 == _T_727 ? _next_reg_T_214 : _GEN_5084; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5181 = 5'h15 == _T_727 ? _next_reg_T_214 : _GEN_5085; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5182 = 5'h16 == _T_727 ? _next_reg_T_214 : _GEN_5086; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5183 = 5'h17 == _T_727 ? _next_reg_T_214 : _GEN_5087; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5184 = 5'h18 == _T_727 ? _next_reg_T_214 : _GEN_5088; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5185 = 5'h19 == _T_727 ? _next_reg_T_214 : _GEN_5089; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5186 = 5'h1a == _T_727 ? _next_reg_T_214 : _GEN_5090; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5187 = 5'h1b == _T_727 ? _next_reg_T_214 : _GEN_5091; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5188 = 5'h1c == _T_727 ? _next_reg_T_214 : _GEN_5092; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5189 = 5'h1d == _T_727 ? _next_reg_T_214 : _GEN_5093; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5190 = 5'h1e == _T_727 ? _next_reg_T_214 : _GEN_5094; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5191 = 5'h1f == _T_727 ? _next_reg_T_214 : _GEN_5095; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_5200 = _T_929 ? _GEN_5161 : _GEN_5065; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5201 = _T_929 ? _GEN_5162 : _GEN_5066; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5202 = _T_929 ? _GEN_5163 : _GEN_5067; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5203 = _T_929 ? _GEN_5164 : _GEN_5068; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5204 = _T_929 ? _GEN_5165 : _GEN_5069; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5205 = _T_929 ? _GEN_5166 : _GEN_5070; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5206 = _T_929 ? _GEN_5167 : _GEN_5071; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5207 = _T_929 ? _GEN_5168 : _GEN_5072; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5208 = _T_929 ? _GEN_5169 : _GEN_5073; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5209 = _T_929 ? _GEN_5170 : _GEN_5074; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5210 = _T_929 ? _GEN_5171 : _GEN_5075; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5211 = _T_929 ? _GEN_5172 : _GEN_5076; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5212 = _T_929 ? _GEN_5173 : _GEN_5077; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5213 = _T_929 ? _GEN_5174 : _GEN_5078; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5214 = _T_929 ? _GEN_5175 : _GEN_5079; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5215 = _T_929 ? _GEN_5176 : _GEN_5080; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5216 = _T_929 ? _GEN_5177 : _GEN_5081; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5217 = _T_929 ? _GEN_5178 : _GEN_5082; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5218 = _T_929 ? _GEN_5179 : _GEN_5083; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5219 = _T_929 ? _GEN_5180 : _GEN_5084; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5220 = _T_929 ? _GEN_5181 : _GEN_5085; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5221 = _T_929 ? _GEN_5182 : _GEN_5086; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5222 = _T_929 ? _GEN_5183 : _GEN_5087; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5223 = _T_929 ? _GEN_5184 : _GEN_5088; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5224 = _T_929 ? _GEN_5185 : _GEN_5089; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5225 = _T_929 ? _GEN_5186 : _GEN_5090; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5226 = _T_929 ? _GEN_5187 : _GEN_5091; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5227 = _T_929 ? _GEN_5188 : _GEN_5092; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5228 = _T_929 ? _GEN_5189 : _GEN_5093; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5229 = _T_929 ? _GEN_5190 : _GEN_5094; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_5230 = _T_929 ? _GEN_5191 : _GEN_5095; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _next_reg_T_217 = _GEN_4675 | _GEN_4116; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:79]
  wire [63:0] _GEN_5296 = 5'h1 == _T_727 ? _next_reg_T_217 : _GEN_5200; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5297 = 5'h2 == _T_727 ? _next_reg_T_217 : _GEN_5201; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5298 = 5'h3 == _T_727 ? _next_reg_T_217 : _GEN_5202; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5299 = 5'h4 == _T_727 ? _next_reg_T_217 : _GEN_5203; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5300 = 5'h5 == _T_727 ? _next_reg_T_217 : _GEN_5204; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5301 = 5'h6 == _T_727 ? _next_reg_T_217 : _GEN_5205; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5302 = 5'h7 == _T_727 ? _next_reg_T_217 : _GEN_5206; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5303 = 5'h8 == _T_727 ? _next_reg_T_217 : _GEN_5207; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5304 = 5'h9 == _T_727 ? _next_reg_T_217 : _GEN_5208; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5305 = 5'ha == _T_727 ? _next_reg_T_217 : _GEN_5209; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5306 = 5'hb == _T_727 ? _next_reg_T_217 : _GEN_5210; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5307 = 5'hc == _T_727 ? _next_reg_T_217 : _GEN_5211; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5308 = 5'hd == _T_727 ? _next_reg_T_217 : _GEN_5212; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5309 = 5'he == _T_727 ? _next_reg_T_217 : _GEN_5213; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5310 = 5'hf == _T_727 ? _next_reg_T_217 : _GEN_5214; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5311 = 5'h10 == _T_727 ? _next_reg_T_217 : _GEN_5215; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5312 = 5'h11 == _T_727 ? _next_reg_T_217 : _GEN_5216; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5313 = 5'h12 == _T_727 ? _next_reg_T_217 : _GEN_5217; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5314 = 5'h13 == _T_727 ? _next_reg_T_217 : _GEN_5218; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5315 = 5'h14 == _T_727 ? _next_reg_T_217 : _GEN_5219; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5316 = 5'h15 == _T_727 ? _next_reg_T_217 : _GEN_5220; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5317 = 5'h16 == _T_727 ? _next_reg_T_217 : _GEN_5221; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5318 = 5'h17 == _T_727 ? _next_reg_T_217 : _GEN_5222; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5319 = 5'h18 == _T_727 ? _next_reg_T_217 : _GEN_5223; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5320 = 5'h19 == _T_727 ? _next_reg_T_217 : _GEN_5224; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5321 = 5'h1a == _T_727 ? _next_reg_T_217 : _GEN_5225; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5322 = 5'h1b == _T_727 ? _next_reg_T_217 : _GEN_5226; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5323 = 5'h1c == _T_727 ? _next_reg_T_217 : _GEN_5227; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5324 = 5'h1d == _T_727 ? _next_reg_T_217 : _GEN_5228; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5325 = 5'h1e == _T_727 ? _next_reg_T_217 : _GEN_5229; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5326 = 5'h1f == _T_727 ? _next_reg_T_217 : _GEN_5230; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_5335 = _T_937 ? _GEN_5296 : _GEN_5200; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5336 = _T_937 ? _GEN_5297 : _GEN_5201; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5337 = _T_937 ? _GEN_5298 : _GEN_5202; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5338 = _T_937 ? _GEN_5299 : _GEN_5203; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5339 = _T_937 ? _GEN_5300 : _GEN_5204; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5340 = _T_937 ? _GEN_5301 : _GEN_5205; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5341 = _T_937 ? _GEN_5302 : _GEN_5206; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5342 = _T_937 ? _GEN_5303 : _GEN_5207; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5343 = _T_937 ? _GEN_5304 : _GEN_5208; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5344 = _T_937 ? _GEN_5305 : _GEN_5209; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5345 = _T_937 ? _GEN_5306 : _GEN_5210; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5346 = _T_937 ? _GEN_5307 : _GEN_5211; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5347 = _T_937 ? _GEN_5308 : _GEN_5212; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5348 = _T_937 ? _GEN_5309 : _GEN_5213; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5349 = _T_937 ? _GEN_5310 : _GEN_5214; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5350 = _T_937 ? _GEN_5311 : _GEN_5215; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5351 = _T_937 ? _GEN_5312 : _GEN_5216; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5352 = _T_937 ? _GEN_5313 : _GEN_5217; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5353 = _T_937 ? _GEN_5314 : _GEN_5218; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5354 = _T_937 ? _GEN_5315 : _GEN_5219; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5355 = _T_937 ? _GEN_5316 : _GEN_5220; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5356 = _T_937 ? _GEN_5317 : _GEN_5221; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5357 = _T_937 ? _GEN_5318 : _GEN_5222; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5358 = _T_937 ? _GEN_5319 : _GEN_5223; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5359 = _T_937 ? _GEN_5320 : _GEN_5224; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5360 = _T_937 ? _GEN_5321 : _GEN_5225; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5361 = _T_937 ? _GEN_5322 : _GEN_5226; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5362 = _T_937 ? _GEN_5323 : _GEN_5227; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5363 = _T_937 ? _GEN_5324 : _GEN_5228; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5364 = _T_937 ? _GEN_5325 : _GEN_5229; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_5365 = _T_937 ? _GEN_5326 : _GEN_5230; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _next_reg_T_220 = _GEN_4675 ^ _GEN_4116; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:79]
  wire [63:0] _GEN_5431 = 5'h1 == _T_727 ? _next_reg_T_220 : _GEN_5335; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5432 = 5'h2 == _T_727 ? _next_reg_T_220 : _GEN_5336; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5433 = 5'h3 == _T_727 ? _next_reg_T_220 : _GEN_5337; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5434 = 5'h4 == _T_727 ? _next_reg_T_220 : _GEN_5338; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5435 = 5'h5 == _T_727 ? _next_reg_T_220 : _GEN_5339; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5436 = 5'h6 == _T_727 ? _next_reg_T_220 : _GEN_5340; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5437 = 5'h7 == _T_727 ? _next_reg_T_220 : _GEN_5341; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5438 = 5'h8 == _T_727 ? _next_reg_T_220 : _GEN_5342; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5439 = 5'h9 == _T_727 ? _next_reg_T_220 : _GEN_5343; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5440 = 5'ha == _T_727 ? _next_reg_T_220 : _GEN_5344; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5441 = 5'hb == _T_727 ? _next_reg_T_220 : _GEN_5345; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5442 = 5'hc == _T_727 ? _next_reg_T_220 : _GEN_5346; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5443 = 5'hd == _T_727 ? _next_reg_T_220 : _GEN_5347; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5444 = 5'he == _T_727 ? _next_reg_T_220 : _GEN_5348; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5445 = 5'hf == _T_727 ? _next_reg_T_220 : _GEN_5349; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5446 = 5'h10 == _T_727 ? _next_reg_T_220 : _GEN_5350; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5447 = 5'h11 == _T_727 ? _next_reg_T_220 : _GEN_5351; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5448 = 5'h12 == _T_727 ? _next_reg_T_220 : _GEN_5352; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5449 = 5'h13 == _T_727 ? _next_reg_T_220 : _GEN_5353; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5450 = 5'h14 == _T_727 ? _next_reg_T_220 : _GEN_5354; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5451 = 5'h15 == _T_727 ? _next_reg_T_220 : _GEN_5355; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5452 = 5'h16 == _T_727 ? _next_reg_T_220 : _GEN_5356; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5453 = 5'h17 == _T_727 ? _next_reg_T_220 : _GEN_5357; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5454 = 5'h18 == _T_727 ? _next_reg_T_220 : _GEN_5358; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5455 = 5'h19 == _T_727 ? _next_reg_T_220 : _GEN_5359; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5456 = 5'h1a == _T_727 ? _next_reg_T_220 : _GEN_5360; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5457 = 5'h1b == _T_727 ? _next_reg_T_220 : _GEN_5361; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5458 = 5'h1c == _T_727 ? _next_reg_T_220 : _GEN_5362; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5459 = 5'h1d == _T_727 ? _next_reg_T_220 : _GEN_5363; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5460 = 5'h1e == _T_727 ? _next_reg_T_220 : _GEN_5364; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5461 = 5'h1f == _T_727 ? _next_reg_T_220 : _GEN_5365; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_5470 = _T_945 ? _GEN_5431 : _GEN_5335; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5471 = _T_945 ? _GEN_5432 : _GEN_5336; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5472 = _T_945 ? _GEN_5433 : _GEN_5337; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5473 = _T_945 ? _GEN_5434 : _GEN_5338; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5474 = _T_945 ? _GEN_5435 : _GEN_5339; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5475 = _T_945 ? _GEN_5436 : _GEN_5340; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5476 = _T_945 ? _GEN_5437 : _GEN_5341; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5477 = _T_945 ? _GEN_5438 : _GEN_5342; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5478 = _T_945 ? _GEN_5439 : _GEN_5343; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5479 = _T_945 ? _GEN_5440 : _GEN_5344; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5480 = _T_945 ? _GEN_5441 : _GEN_5345; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5481 = _T_945 ? _GEN_5442 : _GEN_5346; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5482 = _T_945 ? _GEN_5443 : _GEN_5347; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5483 = _T_945 ? _GEN_5444 : _GEN_5348; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5484 = _T_945 ? _GEN_5445 : _GEN_5349; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5485 = _T_945 ? _GEN_5446 : _GEN_5350; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5486 = _T_945 ? _GEN_5447 : _GEN_5351; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5487 = _T_945 ? _GEN_5448 : _GEN_5352; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5488 = _T_945 ? _GEN_5449 : _GEN_5353; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5489 = _T_945 ? _GEN_5450 : _GEN_5354; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5490 = _T_945 ? _GEN_5451 : _GEN_5355; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5491 = _T_945 ? _GEN_5452 : _GEN_5356; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5492 = _T_945 ? _GEN_5453 : _GEN_5357; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5493 = _T_945 ? _GEN_5454 : _GEN_5358; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5494 = _T_945 ? _GEN_5455 : _GEN_5359; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5495 = _T_945 ? _GEN_5456 : _GEN_5360; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5496 = _T_945 ? _GEN_5457 : _GEN_5361; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5497 = _T_945 ? _GEN_5458 : _GEN_5362; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5498 = _T_945 ? _GEN_5459 : _GEN_5363; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5499 = _T_945 ? _GEN_5460 : _GEN_5364; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_5500 = _T_945 ? _GEN_5461 : _GEN_5365; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _next_reg_T_224 = _GEN_4675 - _GEN_4116; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:79]
  wire [63:0] _GEN_5566 = 5'h1 == _T_727 ? _next_reg_T_224 : _GEN_5470; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5567 = 5'h2 == _T_727 ? _next_reg_T_224 : _GEN_5471; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5568 = 5'h3 == _T_727 ? _next_reg_T_224 : _GEN_5472; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5569 = 5'h4 == _T_727 ? _next_reg_T_224 : _GEN_5473; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5570 = 5'h5 == _T_727 ? _next_reg_T_224 : _GEN_5474; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5571 = 5'h6 == _T_727 ? _next_reg_T_224 : _GEN_5475; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5572 = 5'h7 == _T_727 ? _next_reg_T_224 : _GEN_5476; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5573 = 5'h8 == _T_727 ? _next_reg_T_224 : _GEN_5477; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5574 = 5'h9 == _T_727 ? _next_reg_T_224 : _GEN_5478; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5575 = 5'ha == _T_727 ? _next_reg_T_224 : _GEN_5479; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5576 = 5'hb == _T_727 ? _next_reg_T_224 : _GEN_5480; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5577 = 5'hc == _T_727 ? _next_reg_T_224 : _GEN_5481; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5578 = 5'hd == _T_727 ? _next_reg_T_224 : _GEN_5482; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5579 = 5'he == _T_727 ? _next_reg_T_224 : _GEN_5483; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5580 = 5'hf == _T_727 ? _next_reg_T_224 : _GEN_5484; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5581 = 5'h10 == _T_727 ? _next_reg_T_224 : _GEN_5485; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5582 = 5'h11 == _T_727 ? _next_reg_T_224 : _GEN_5486; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5583 = 5'h12 == _T_727 ? _next_reg_T_224 : _GEN_5487; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5584 = 5'h13 == _T_727 ? _next_reg_T_224 : _GEN_5488; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5585 = 5'h14 == _T_727 ? _next_reg_T_224 : _GEN_5489; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5586 = 5'h15 == _T_727 ? _next_reg_T_224 : _GEN_5490; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5587 = 5'h16 == _T_727 ? _next_reg_T_224 : _GEN_5491; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5588 = 5'h17 == _T_727 ? _next_reg_T_224 : _GEN_5492; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5589 = 5'h18 == _T_727 ? _next_reg_T_224 : _GEN_5493; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5590 = 5'h19 == _T_727 ? _next_reg_T_224 : _GEN_5494; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5591 = 5'h1a == _T_727 ? _next_reg_T_224 : _GEN_5495; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5592 = 5'h1b == _T_727 ? _next_reg_T_224 : _GEN_5496; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5593 = 5'h1c == _T_727 ? _next_reg_T_224 : _GEN_5497; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5594 = 5'h1d == _T_727 ? _next_reg_T_224 : _GEN_5498; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5595 = 5'h1e == _T_727 ? _next_reg_T_224 : _GEN_5499; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5596 = 5'h1f == _T_727 ? _next_reg_T_224 : _GEN_5500; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_5605 = _T_953 ? _GEN_5566 : _GEN_5470; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5606 = _T_953 ? _GEN_5567 : _GEN_5471; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5607 = _T_953 ? _GEN_5568 : _GEN_5472; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5608 = _T_953 ? _GEN_5569 : _GEN_5473; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5609 = _T_953 ? _GEN_5570 : _GEN_5474; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5610 = _T_953 ? _GEN_5571 : _GEN_5475; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5611 = _T_953 ? _GEN_5572 : _GEN_5476; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5612 = _T_953 ? _GEN_5573 : _GEN_5477; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5613 = _T_953 ? _GEN_5574 : _GEN_5478; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5614 = _T_953 ? _GEN_5575 : _GEN_5479; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5615 = _T_953 ? _GEN_5576 : _GEN_5480; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5616 = _T_953 ? _GEN_5577 : _GEN_5481; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5617 = _T_953 ? _GEN_5578 : _GEN_5482; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5618 = _T_953 ? _GEN_5579 : _GEN_5483; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5619 = _T_953 ? _GEN_5580 : _GEN_5484; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5620 = _T_953 ? _GEN_5581 : _GEN_5485; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5621 = _T_953 ? _GEN_5582 : _GEN_5486; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5622 = _T_953 ? _GEN_5583 : _GEN_5487; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5623 = _T_953 ? _GEN_5584 : _GEN_5488; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5624 = _T_953 ? _GEN_5585 : _GEN_5489; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5625 = _T_953 ? _GEN_5586 : _GEN_5490; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5626 = _T_953 ? _GEN_5587 : _GEN_5491; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5627 = _T_953 ? _GEN_5588 : _GEN_5492; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5628 = _T_953 ? _GEN_5589 : _GEN_5493; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5629 = _T_953 ? _GEN_5590 : _GEN_5494; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5630 = _T_953 ? _GEN_5591 : _GEN_5495; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5631 = _T_953 ? _GEN_5592 : _GEN_5496; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5632 = _T_953 ? _GEN_5593 : _GEN_5497; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5633 = _T_953 ? _GEN_5594 : _GEN_5498; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5634 = _T_953 ? _GEN_5595 : _GEN_5499; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5635 = _T_953 ? _GEN_5596 : _GEN_5500; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_5644 = 5'h1 == rd ? _next_reg_T_177 : _GEN_5605; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5645 = 5'h2 == rd ? _next_reg_T_177 : _GEN_5606; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5646 = 5'h3 == rd ? _next_reg_T_177 : _GEN_5607; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5647 = 5'h4 == rd ? _next_reg_T_177 : _GEN_5608; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5648 = 5'h5 == rd ? _next_reg_T_177 : _GEN_5609; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5649 = 5'h6 == rd ? _next_reg_T_177 : _GEN_5610; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5650 = 5'h7 == rd ? _next_reg_T_177 : _GEN_5611; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5651 = 5'h8 == rd ? _next_reg_T_177 : _GEN_5612; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5652 = 5'h9 == rd ? _next_reg_T_177 : _GEN_5613; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5653 = 5'ha == rd ? _next_reg_T_177 : _GEN_5614; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5654 = 5'hb == rd ? _next_reg_T_177 : _GEN_5615; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5655 = 5'hc == rd ? _next_reg_T_177 : _GEN_5616; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5656 = 5'hd == rd ? _next_reg_T_177 : _GEN_5617; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5657 = 5'he == rd ? _next_reg_T_177 : _GEN_5618; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5658 = 5'hf == rd ? _next_reg_T_177 : _GEN_5619; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5659 = 5'h10 == rd ? _next_reg_T_177 : _GEN_5620; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5660 = 5'h11 == rd ? _next_reg_T_177 : _GEN_5621; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5661 = 5'h12 == rd ? _next_reg_T_177 : _GEN_5622; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5662 = 5'h13 == rd ? _next_reg_T_177 : _GEN_5623; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5663 = 5'h14 == rd ? _next_reg_T_177 : _GEN_5624; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5664 = 5'h15 == rd ? _next_reg_T_177 : _GEN_5625; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5665 = 5'h16 == rd ? _next_reg_T_177 : _GEN_5626; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5666 = 5'h17 == rd ? _next_reg_T_177 : _GEN_5627; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5667 = 5'h18 == rd ? _next_reg_T_177 : _GEN_5628; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5668 = 5'h19 == rd ? _next_reg_T_177 : _GEN_5629; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5669 = 5'h1a == rd ? _next_reg_T_177 : _GEN_5630; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5670 = 5'h1b == rd ? _next_reg_T_177 : _GEN_5631; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5671 = 5'h1c == rd ? _next_reg_T_177 : _GEN_5632; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5672 = 5'h1d == rd ? _next_reg_T_177 : _GEN_5633; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5673 = 5'h1e == rd ? _next_reg_T_177 : _GEN_5634; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_5674 = 5'h1f == rd ? _next_reg_T_177 : _GEN_5635; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire  _GEN_5683 = _T_971 | _GEN_4018; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [63:0] _GEN_5684 = _T_971 ? _next_reg_T_176 : _GEN_4019; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [6:0] _GEN_5685 = _T_971 ? 7'h40 : _GEN_4020; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [63:0] _GEN_5687 = _T_971 ? _GEN_5644 : _GEN_5605; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5688 = _T_971 ? _GEN_5645 : _GEN_5606; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5689 = _T_971 ? _GEN_5646 : _GEN_5607; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5690 = _T_971 ? _GEN_5647 : _GEN_5608; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5691 = _T_971 ? _GEN_5648 : _GEN_5609; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5692 = _T_971 ? _GEN_5649 : _GEN_5610; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5693 = _T_971 ? _GEN_5650 : _GEN_5611; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5694 = _T_971 ? _GEN_5651 : _GEN_5612; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5695 = _T_971 ? _GEN_5652 : _GEN_5613; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5696 = _T_971 ? _GEN_5653 : _GEN_5614; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5697 = _T_971 ? _GEN_5654 : _GEN_5615; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5698 = _T_971 ? _GEN_5655 : _GEN_5616; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5699 = _T_971 ? _GEN_5656 : _GEN_5617; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5700 = _T_971 ? _GEN_5657 : _GEN_5618; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5701 = _T_971 ? _GEN_5658 : _GEN_5619; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5702 = _T_971 ? _GEN_5659 : _GEN_5620; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5703 = _T_971 ? _GEN_5660 : _GEN_5621; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5704 = _T_971 ? _GEN_5661 : _GEN_5622; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5705 = _T_971 ? _GEN_5662 : _GEN_5623; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5706 = _T_971 ? _GEN_5663 : _GEN_5624; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5707 = _T_971 ? _GEN_5664 : _GEN_5625; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5708 = _T_971 ? _GEN_5665 : _GEN_5626; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5709 = _T_971 ? _GEN_5666 : _GEN_5627; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5710 = _T_971 ? _GEN_5667 : _GEN_5628; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5711 = _T_971 ? _GEN_5668 : _GEN_5629; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5712 = _T_971 ? _GEN_5669 : _GEN_5630; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5713 = _T_971 ? _GEN_5670 : _GEN_5631; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5714 = _T_971 ? _GEN_5671 : _GEN_5632; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5715 = _T_971 ? _GEN_5672 : _GEN_5633; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5716 = _T_971 ? _GEN_5673 : _GEN_5634; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_5717 = _T_971 ? _GEN_5674 : _GEN_5635; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire  _GEN_5724 = _T_978 | _GEN_4125; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 82:26]
  wire [63:0] _GEN_5725 = _T_978 ? _next_reg_T_176 : _GEN_4126; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 83:26]
  wire [6:0] _GEN_5726 = _T_978 ? 7'h40 : _GEN_4127; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 84:26]
  wire [63:0] _GEN_5727 = _T_978 ? _GEN_840 : _GEN_4128; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:26]
  wire [63:0] _GEN_5761 = 5'h1 == _T_727 ? _next_reg_T_186 : _GEN_5687; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5762 = 5'h2 == _T_727 ? _next_reg_T_186 : _GEN_5688; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5763 = 5'h3 == _T_727 ? _next_reg_T_186 : _GEN_5689; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5764 = 5'h4 == _T_727 ? _next_reg_T_186 : _GEN_5690; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5765 = 5'h5 == _T_727 ? _next_reg_T_186 : _GEN_5691; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5766 = 5'h6 == _T_727 ? _next_reg_T_186 : _GEN_5692; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5767 = 5'h7 == _T_727 ? _next_reg_T_186 : _GEN_5693; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5768 = 5'h8 == _T_727 ? _next_reg_T_186 : _GEN_5694; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5769 = 5'h9 == _T_727 ? _next_reg_T_186 : _GEN_5695; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5770 = 5'ha == _T_727 ? _next_reg_T_186 : _GEN_5696; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5771 = 5'hb == _T_727 ? _next_reg_T_186 : _GEN_5697; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5772 = 5'hc == _T_727 ? _next_reg_T_186 : _GEN_5698; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5773 = 5'hd == _T_727 ? _next_reg_T_186 : _GEN_5699; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5774 = 5'he == _T_727 ? _next_reg_T_186 : _GEN_5700; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5775 = 5'hf == _T_727 ? _next_reg_T_186 : _GEN_5701; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5776 = 5'h10 == _T_727 ? _next_reg_T_186 : _GEN_5702; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5777 = 5'h11 == _T_727 ? _next_reg_T_186 : _GEN_5703; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5778 = 5'h12 == _T_727 ? _next_reg_T_186 : _GEN_5704; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5779 = 5'h13 == _T_727 ? _next_reg_T_186 : _GEN_5705; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5780 = 5'h14 == _T_727 ? _next_reg_T_186 : _GEN_5706; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5781 = 5'h15 == _T_727 ? _next_reg_T_186 : _GEN_5707; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5782 = 5'h16 == _T_727 ? _next_reg_T_186 : _GEN_5708; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5783 = 5'h17 == _T_727 ? _next_reg_T_186 : _GEN_5709; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5784 = 5'h18 == _T_727 ? _next_reg_T_186 : _GEN_5710; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5785 = 5'h19 == _T_727 ? _next_reg_T_186 : _GEN_5711; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5786 = 5'h1a == _T_727 ? _next_reg_T_186 : _GEN_5712; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5787 = 5'h1b == _T_727 ? _next_reg_T_186 : _GEN_5713; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5788 = 5'h1c == _T_727 ? _next_reg_T_186 : _GEN_5714; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5789 = 5'h1d == _T_727 ? _next_reg_T_186 : _GEN_5715; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5790 = 5'h1e == _T_727 ? _next_reg_T_186 : _GEN_5716; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_5791 = 5'h1f == _T_727 ? _next_reg_T_186 : _GEN_5717; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire  _GEN_5800 = _T_987 | _GEN_5683; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 52:25]
  wire [63:0] _GEN_5801 = _T_987 ? _next_reg_T_185 : _GEN_5684; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 53:25]
  wire [6:0] _GEN_5802 = _T_987 ? 7'h40 : _GEN_5685; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 54:25]
  wire [63:0] _GEN_5804 = _T_987 ? _GEN_5761 : _GEN_5687; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5805 = _T_987 ? _GEN_5762 : _GEN_5688; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5806 = _T_987 ? _GEN_5763 : _GEN_5689; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5807 = _T_987 ? _GEN_5764 : _GEN_5690; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5808 = _T_987 ? _GEN_5765 : _GEN_5691; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5809 = _T_987 ? _GEN_5766 : _GEN_5692; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5810 = _T_987 ? _GEN_5767 : _GEN_5693; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5811 = _T_987 ? _GEN_5768 : _GEN_5694; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5812 = _T_987 ? _GEN_5769 : _GEN_5695; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5813 = _T_987 ? _GEN_5770 : _GEN_5696; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5814 = _T_987 ? _GEN_5771 : _GEN_5697; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5815 = _T_987 ? _GEN_5772 : _GEN_5698; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5816 = _T_987 ? _GEN_5773 : _GEN_5699; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5817 = _T_987 ? _GEN_5774 : _GEN_5700; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5818 = _T_987 ? _GEN_5775 : _GEN_5701; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5819 = _T_987 ? _GEN_5776 : _GEN_5702; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5820 = _T_987 ? _GEN_5777 : _GEN_5703; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5821 = _T_987 ? _GEN_5778 : _GEN_5704; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5822 = _T_987 ? _GEN_5779 : _GEN_5705; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5823 = _T_987 ? _GEN_5780 : _GEN_5706; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5824 = _T_987 ? _GEN_5781 : _GEN_5707; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5825 = _T_987 ? _GEN_5782 : _GEN_5708; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5826 = _T_987 ? _GEN_5783 : _GEN_5709; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5827 = _T_987 ? _GEN_5784 : _GEN_5710; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5828 = _T_987 ? _GEN_5785 : _GEN_5711; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5829 = _T_987 ? _GEN_5786 : _GEN_5712; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5830 = _T_987 ? _GEN_5787 : _GEN_5713; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5831 = _T_987 ? _GEN_5788 : _GEN_5714; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5832 = _T_987 ? _GEN_5789 : _GEN_5715; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5833 = _T_987 ? _GEN_5790 : _GEN_5716; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_5834 = _T_987 ? _GEN_5791 : _GEN_5717; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire  _GEN_5907 = _T_996 | _GEN_5724; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 82:26]
  wire [63:0] _GEN_5908 = _T_996 ? _next_reg_T_185 : _GEN_5725; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 83:26]
  wire [6:0] _GEN_5909 = _T_996 ? 7'h40 : _GEN_5726; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 84:26]
  wire [63:0] _GEN_5910 = _T_996 ? _GEN_4116 : _GEN_5727; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 85:26]
  wire [63:0] _next_reg_T_239 = _GEN_4423 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:44]
  wire  next_reg_signBit_17 = _next_reg_T_239[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_242 = next_reg_signBit_17 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_243 = {_next_reg_T_242,_next_reg_T_239[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_5912 = 5'h1 == rd ? _next_reg_T_243 : _GEN_5804; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5913 = 5'h2 == rd ? _next_reg_T_243 : _GEN_5805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5914 = 5'h3 == rd ? _next_reg_T_243 : _GEN_5806; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5915 = 5'h4 == rd ? _next_reg_T_243 : _GEN_5807; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5916 = 5'h5 == rd ? _next_reg_T_243 : _GEN_5808; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5917 = 5'h6 == rd ? _next_reg_T_243 : _GEN_5809; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5918 = 5'h7 == rd ? _next_reg_T_243 : _GEN_5810; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5919 = 5'h8 == rd ? _next_reg_T_243 : _GEN_5811; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5920 = 5'h9 == rd ? _next_reg_T_243 : _GEN_5812; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5921 = 5'ha == rd ? _next_reg_T_243 : _GEN_5813; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5922 = 5'hb == rd ? _next_reg_T_243 : _GEN_5814; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5923 = 5'hc == rd ? _next_reg_T_243 : _GEN_5815; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5924 = 5'hd == rd ? _next_reg_T_243 : _GEN_5816; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5925 = 5'he == rd ? _next_reg_T_243 : _GEN_5817; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5926 = 5'hf == rd ? _next_reg_T_243 : _GEN_5818; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5927 = 5'h10 == rd ? _next_reg_T_243 : _GEN_5819; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5928 = 5'h11 == rd ? _next_reg_T_243 : _GEN_5820; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5929 = 5'h12 == rd ? _next_reg_T_243 : _GEN_5821; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5930 = 5'h13 == rd ? _next_reg_T_243 : _GEN_5822; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5931 = 5'h14 == rd ? _next_reg_T_243 : _GEN_5823; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5932 = 5'h15 == rd ? _next_reg_T_243 : _GEN_5824; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5933 = 5'h16 == rd ? _next_reg_T_243 : _GEN_5825; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5934 = 5'h17 == rd ? _next_reg_T_243 : _GEN_5826; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5935 = 5'h18 == rd ? _next_reg_T_243 : _GEN_5827; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5936 = 5'h19 == rd ? _next_reg_T_243 : _GEN_5828; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5937 = 5'h1a == rd ? _next_reg_T_243 : _GEN_5829; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5938 = 5'h1b == rd ? _next_reg_T_243 : _GEN_5830; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5939 = 5'h1c == rd ? _next_reg_T_243 : _GEN_5831; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5940 = 5'h1d == rd ? _next_reg_T_243 : _GEN_5832; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5941 = 5'h1e == rd ? _next_reg_T_243 : _GEN_5833; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5942 = 5'h1f == rd ? _next_reg_T_243 : _GEN_5834; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_5952 = _T_1011 ? _GEN_5912 : _GEN_5804; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5953 = _T_1011 ? _GEN_5913 : _GEN_5805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5954 = _T_1011 ? _GEN_5914 : _GEN_5806; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5955 = _T_1011 ? _GEN_5915 : _GEN_5807; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5956 = _T_1011 ? _GEN_5916 : _GEN_5808; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5957 = _T_1011 ? _GEN_5917 : _GEN_5809; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5958 = _T_1011 ? _GEN_5918 : _GEN_5810; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5959 = _T_1011 ? _GEN_5919 : _GEN_5811; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5960 = _T_1011 ? _GEN_5920 : _GEN_5812; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5961 = _T_1011 ? _GEN_5921 : _GEN_5813; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5962 = _T_1011 ? _GEN_5922 : _GEN_5814; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5963 = _T_1011 ? _GEN_5923 : _GEN_5815; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5964 = _T_1011 ? _GEN_5924 : _GEN_5816; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5965 = _T_1011 ? _GEN_5925 : _GEN_5817; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5966 = _T_1011 ? _GEN_5926 : _GEN_5818; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5967 = _T_1011 ? _GEN_5927 : _GEN_5819; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5968 = _T_1011 ? _GEN_5928 : _GEN_5820; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5969 = _T_1011 ? _GEN_5929 : _GEN_5821; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5970 = _T_1011 ? _GEN_5930 : _GEN_5822; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5971 = _T_1011 ? _GEN_5931 : _GEN_5823; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5972 = _T_1011 ? _GEN_5932 : _GEN_5824; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5973 = _T_1011 ? _GEN_5933 : _GEN_5825; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5974 = _T_1011 ? _GEN_5934 : _GEN_5826; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5975 = _T_1011 ? _GEN_5935 : _GEN_5827; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5976 = _T_1011 ? _GEN_5936 : _GEN_5828; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5977 = _T_1011 ? _GEN_5937 : _GEN_5829; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5978 = _T_1011 ? _GEN_5938 : _GEN_5830; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5979 = _T_1011 ? _GEN_5939 : _GEN_5831; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5980 = _T_1011 ? _GEN_5940 : _GEN_5832; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5981 = _T_1011 ? _GEN_5941 : _GEN_5833; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_5982 = _T_1011 ? _GEN_5942 : _GEN_5834; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [31:0] _next_reg_T_249 = _GEN_4675[31:0] + _GEN_4116[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:66]
  wire  next_reg_signBit_18 = _next_reg_T_249[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_251 = next_reg_signBit_18 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_252 = {_next_reg_T_251,_next_reg_T_249}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_6048 = 5'h1 == _T_727 ? _next_reg_T_252 : _GEN_5952; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6049 = 5'h2 == _T_727 ? _next_reg_T_252 : _GEN_5953; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6050 = 5'h3 == _T_727 ? _next_reg_T_252 : _GEN_5954; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6051 = 5'h4 == _T_727 ? _next_reg_T_252 : _GEN_5955; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6052 = 5'h5 == _T_727 ? _next_reg_T_252 : _GEN_5956; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6053 = 5'h6 == _T_727 ? _next_reg_T_252 : _GEN_5957; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6054 = 5'h7 == _T_727 ? _next_reg_T_252 : _GEN_5958; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6055 = 5'h8 == _T_727 ? _next_reg_T_252 : _GEN_5959; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6056 = 5'h9 == _T_727 ? _next_reg_T_252 : _GEN_5960; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6057 = 5'ha == _T_727 ? _next_reg_T_252 : _GEN_5961; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6058 = 5'hb == _T_727 ? _next_reg_T_252 : _GEN_5962; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6059 = 5'hc == _T_727 ? _next_reg_T_252 : _GEN_5963; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6060 = 5'hd == _T_727 ? _next_reg_T_252 : _GEN_5964; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6061 = 5'he == _T_727 ? _next_reg_T_252 : _GEN_5965; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6062 = 5'hf == _T_727 ? _next_reg_T_252 : _GEN_5966; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6063 = 5'h10 == _T_727 ? _next_reg_T_252 : _GEN_5967; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6064 = 5'h11 == _T_727 ? _next_reg_T_252 : _GEN_5968; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6065 = 5'h12 == _T_727 ? _next_reg_T_252 : _GEN_5969; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6066 = 5'h13 == _T_727 ? _next_reg_T_252 : _GEN_5970; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6067 = 5'h14 == _T_727 ? _next_reg_T_252 : _GEN_5971; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6068 = 5'h15 == _T_727 ? _next_reg_T_252 : _GEN_5972; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6069 = 5'h16 == _T_727 ? _next_reg_T_252 : _GEN_5973; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6070 = 5'h17 == _T_727 ? _next_reg_T_252 : _GEN_5974; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6071 = 5'h18 == _T_727 ? _next_reg_T_252 : _GEN_5975; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6072 = 5'h19 == _T_727 ? _next_reg_T_252 : _GEN_5976; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6073 = 5'h1a == _T_727 ? _next_reg_T_252 : _GEN_5977; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6074 = 5'h1b == _T_727 ? _next_reg_T_252 : _GEN_5978; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6075 = 5'h1c == _T_727 ? _next_reg_T_252 : _GEN_5979; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6076 = 5'h1d == _T_727 ? _next_reg_T_252 : _GEN_5980; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6077 = 5'h1e == _T_727 ? _next_reg_T_252 : _GEN_5981; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6078 = 5'h1f == _T_727 ? _next_reg_T_252 : _GEN_5982; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_6087 = _T_1018 ? _GEN_6048 : _GEN_5952; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6088 = _T_1018 ? _GEN_6049 : _GEN_5953; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6089 = _T_1018 ? _GEN_6050 : _GEN_5954; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6090 = _T_1018 ? _GEN_6051 : _GEN_5955; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6091 = _T_1018 ? _GEN_6052 : _GEN_5956; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6092 = _T_1018 ? _GEN_6053 : _GEN_5957; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6093 = _T_1018 ? _GEN_6054 : _GEN_5958; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6094 = _T_1018 ? _GEN_6055 : _GEN_5959; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6095 = _T_1018 ? _GEN_6056 : _GEN_5960; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6096 = _T_1018 ? _GEN_6057 : _GEN_5961; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6097 = _T_1018 ? _GEN_6058 : _GEN_5962; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6098 = _T_1018 ? _GEN_6059 : _GEN_5963; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6099 = _T_1018 ? _GEN_6060 : _GEN_5964; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6100 = _T_1018 ? _GEN_6061 : _GEN_5965; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6101 = _T_1018 ? _GEN_6062 : _GEN_5966; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6102 = _T_1018 ? _GEN_6063 : _GEN_5967; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6103 = _T_1018 ? _GEN_6064 : _GEN_5968; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6104 = _T_1018 ? _GEN_6065 : _GEN_5969; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6105 = _T_1018 ? _GEN_6066 : _GEN_5970; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6106 = _T_1018 ? _GEN_6067 : _GEN_5971; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6107 = _T_1018 ? _GEN_6068 : _GEN_5972; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6108 = _T_1018 ? _GEN_6069 : _GEN_5973; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6109 = _T_1018 ? _GEN_6070 : _GEN_5974; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6110 = _T_1018 ? _GEN_6071 : _GEN_5975; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6111 = _T_1018 ? _GEN_6072 : _GEN_5976; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6112 = _T_1018 ? _GEN_6073 : _GEN_5977; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6113 = _T_1018 ? _GEN_6074 : _GEN_5978; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6114 = _T_1018 ? _GEN_6075 : _GEN_5979; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6115 = _T_1018 ? _GEN_6076 : _GEN_5980; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6116 = _T_1018 ? _GEN_6077 : _GEN_5981; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_6117 = _T_1018 ? _GEN_6078 : _GEN_5982; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [31:0] _next_reg_T_258 = _GEN_4675[31:0] - _GEN_4116[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:66]
  wire  next_reg_signBit_19 = _next_reg_T_258[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_260 = next_reg_signBit_19 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_261 = {_next_reg_T_260,_next_reg_T_258}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_6183 = 5'h1 == _T_727 ? _next_reg_T_261 : _GEN_6087; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6184 = 5'h2 == _T_727 ? _next_reg_T_261 : _GEN_6088; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6185 = 5'h3 == _T_727 ? _next_reg_T_261 : _GEN_6089; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6186 = 5'h4 == _T_727 ? _next_reg_T_261 : _GEN_6090; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6187 = 5'h5 == _T_727 ? _next_reg_T_261 : _GEN_6091; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6188 = 5'h6 == _T_727 ? _next_reg_T_261 : _GEN_6092; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6189 = 5'h7 == _T_727 ? _next_reg_T_261 : _GEN_6093; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6190 = 5'h8 == _T_727 ? _next_reg_T_261 : _GEN_6094; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6191 = 5'h9 == _T_727 ? _next_reg_T_261 : _GEN_6095; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6192 = 5'ha == _T_727 ? _next_reg_T_261 : _GEN_6096; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6193 = 5'hb == _T_727 ? _next_reg_T_261 : _GEN_6097; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6194 = 5'hc == _T_727 ? _next_reg_T_261 : _GEN_6098; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6195 = 5'hd == _T_727 ? _next_reg_T_261 : _GEN_6099; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6196 = 5'he == _T_727 ? _next_reg_T_261 : _GEN_6100; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6197 = 5'hf == _T_727 ? _next_reg_T_261 : _GEN_6101; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6198 = 5'h10 == _T_727 ? _next_reg_T_261 : _GEN_6102; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6199 = 5'h11 == _T_727 ? _next_reg_T_261 : _GEN_6103; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6200 = 5'h12 == _T_727 ? _next_reg_T_261 : _GEN_6104; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6201 = 5'h13 == _T_727 ? _next_reg_T_261 : _GEN_6105; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6202 = 5'h14 == _T_727 ? _next_reg_T_261 : _GEN_6106; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6203 = 5'h15 == _T_727 ? _next_reg_T_261 : _GEN_6107; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6204 = 5'h16 == _T_727 ? _next_reg_T_261 : _GEN_6108; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6205 = 5'h17 == _T_727 ? _next_reg_T_261 : _GEN_6109; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6206 = 5'h18 == _T_727 ? _next_reg_T_261 : _GEN_6110; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6207 = 5'h19 == _T_727 ? _next_reg_T_261 : _GEN_6111; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6208 = 5'h1a == _T_727 ? _next_reg_T_261 : _GEN_6112; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6209 = 5'h1b == _T_727 ? _next_reg_T_261 : _GEN_6113; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6210 = 5'h1c == _T_727 ? _next_reg_T_261 : _GEN_6114; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6211 = 5'h1d == _T_727 ? _next_reg_T_261 : _GEN_6115; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6212 = 5'h1e == _T_727 ? _next_reg_T_261 : _GEN_6116; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6213 = 5'h1f == _T_727 ? _next_reg_T_261 : _GEN_6117; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_6222 = _T_1026 ? _GEN_6183 : _GEN_6087; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6223 = _T_1026 ? _GEN_6184 : _GEN_6088; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6224 = _T_1026 ? _GEN_6185 : _GEN_6089; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6225 = _T_1026 ? _GEN_6186 : _GEN_6090; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6226 = _T_1026 ? _GEN_6187 : _GEN_6091; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6227 = _T_1026 ? _GEN_6188 : _GEN_6092; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6228 = _T_1026 ? _GEN_6189 : _GEN_6093; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6229 = _T_1026 ? _GEN_6190 : _GEN_6094; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6230 = _T_1026 ? _GEN_6191 : _GEN_6095; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6231 = _T_1026 ? _GEN_6192 : _GEN_6096; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6232 = _T_1026 ? _GEN_6193 : _GEN_6097; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6233 = _T_1026 ? _GEN_6194 : _GEN_6098; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6234 = _T_1026 ? _GEN_6195 : _GEN_6099; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6235 = _T_1026 ? _GEN_6196 : _GEN_6100; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6236 = _T_1026 ? _GEN_6197 : _GEN_6101; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6237 = _T_1026 ? _GEN_6198 : _GEN_6102; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6238 = _T_1026 ? _GEN_6199 : _GEN_6103; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6239 = _T_1026 ? _GEN_6200 : _GEN_6104; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6240 = _T_1026 ? _GEN_6201 : _GEN_6105; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6241 = _T_1026 ? _GEN_6202 : _GEN_6106; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6242 = _T_1026 ? _GEN_6203 : _GEN_6107; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6243 = _T_1026 ? _GEN_6204 : _GEN_6108; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6244 = _T_1026 ? _GEN_6205 : _GEN_6109; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6245 = _T_1026 ? _GEN_6206 : _GEN_6110; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6246 = _T_1026 ? _GEN_6207 : _GEN_6111; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6247 = _T_1026 ? _GEN_6208 : _GEN_6112; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6248 = _T_1026 ? _GEN_6209 : _GEN_6113; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6249 = _T_1026 ? _GEN_6210 : _GEN_6114; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6250 = _T_1026 ? _GEN_6211 : _GEN_6115; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6251 = _T_1026 ? _GEN_6212 : _GEN_6116; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_6252 = _T_1026 ? _GEN_6213 : _GEN_6117; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [127:0] _next_reg_T_262 = _GEN_31 * _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:65]
  wire [63:0] _GEN_6254 = 5'h1 == rd ? _next_reg_T_262[63:0] : _GEN_6222; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6255 = 5'h2 == rd ? _next_reg_T_262[63:0] : _GEN_6223; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6256 = 5'h3 == rd ? _next_reg_T_262[63:0] : _GEN_6224; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6257 = 5'h4 == rd ? _next_reg_T_262[63:0] : _GEN_6225; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6258 = 5'h5 == rd ? _next_reg_T_262[63:0] : _GEN_6226; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6259 = 5'h6 == rd ? _next_reg_T_262[63:0] : _GEN_6227; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6260 = 5'h7 == rd ? _next_reg_T_262[63:0] : _GEN_6228; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6261 = 5'h8 == rd ? _next_reg_T_262[63:0] : _GEN_6229; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6262 = 5'h9 == rd ? _next_reg_T_262[63:0] : _GEN_6230; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6263 = 5'ha == rd ? _next_reg_T_262[63:0] : _GEN_6231; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6264 = 5'hb == rd ? _next_reg_T_262[63:0] : _GEN_6232; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6265 = 5'hc == rd ? _next_reg_T_262[63:0] : _GEN_6233; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6266 = 5'hd == rd ? _next_reg_T_262[63:0] : _GEN_6234; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6267 = 5'he == rd ? _next_reg_T_262[63:0] : _GEN_6235; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6268 = 5'hf == rd ? _next_reg_T_262[63:0] : _GEN_6236; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6269 = 5'h10 == rd ? _next_reg_T_262[63:0] : _GEN_6237; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6270 = 5'h11 == rd ? _next_reg_T_262[63:0] : _GEN_6238; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6271 = 5'h12 == rd ? _next_reg_T_262[63:0] : _GEN_6239; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6272 = 5'h13 == rd ? _next_reg_T_262[63:0] : _GEN_6240; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6273 = 5'h14 == rd ? _next_reg_T_262[63:0] : _GEN_6241; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6274 = 5'h15 == rd ? _next_reg_T_262[63:0] : _GEN_6242; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6275 = 5'h16 == rd ? _next_reg_T_262[63:0] : _GEN_6243; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6276 = 5'h17 == rd ? _next_reg_T_262[63:0] : _GEN_6244; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6277 = 5'h18 == rd ? _next_reg_T_262[63:0] : _GEN_6245; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6278 = 5'h19 == rd ? _next_reg_T_262[63:0] : _GEN_6246; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6279 = 5'h1a == rd ? _next_reg_T_262[63:0] : _GEN_6247; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6280 = 5'h1b == rd ? _next_reg_T_262[63:0] : _GEN_6248; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6281 = 5'h1c == rd ? _next_reg_T_262[63:0] : _GEN_6249; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6282 = 5'h1d == rd ? _next_reg_T_262[63:0] : _GEN_6250; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6283 = 5'h1e == rd ? _next_reg_T_262[63:0] : _GEN_6251; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6284 = 5'h1f == rd ? _next_reg_T_262[63:0] : _GEN_6252; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_6293 = _T_1034 ? _GEN_6254 : _GEN_6222; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6294 = _T_1034 ? _GEN_6255 : _GEN_6223; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6295 = _T_1034 ? _GEN_6256 : _GEN_6224; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6296 = _T_1034 ? _GEN_6257 : _GEN_6225; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6297 = _T_1034 ? _GEN_6258 : _GEN_6226; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6298 = _T_1034 ? _GEN_6259 : _GEN_6227; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6299 = _T_1034 ? _GEN_6260 : _GEN_6228; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6300 = _T_1034 ? _GEN_6261 : _GEN_6229; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6301 = _T_1034 ? _GEN_6262 : _GEN_6230; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6302 = _T_1034 ? _GEN_6263 : _GEN_6231; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6303 = _T_1034 ? _GEN_6264 : _GEN_6232; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6304 = _T_1034 ? _GEN_6265 : _GEN_6233; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6305 = _T_1034 ? _GEN_6266 : _GEN_6234; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6306 = _T_1034 ? _GEN_6267 : _GEN_6235; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6307 = _T_1034 ? _GEN_6268 : _GEN_6236; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6308 = _T_1034 ? _GEN_6269 : _GEN_6237; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6309 = _T_1034 ? _GEN_6270 : _GEN_6238; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6310 = _T_1034 ? _GEN_6271 : _GEN_6239; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6311 = _T_1034 ? _GEN_6272 : _GEN_6240; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6312 = _T_1034 ? _GEN_6273 : _GEN_6241; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6313 = _T_1034 ? _GEN_6274 : _GEN_6242; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6314 = _T_1034 ? _GEN_6275 : _GEN_6243; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6315 = _T_1034 ? _GEN_6276 : _GEN_6244; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6316 = _T_1034 ? _GEN_6277 : _GEN_6245; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6317 = _T_1034 ? _GEN_6278 : _GEN_6246; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6318 = _T_1034 ? _GEN_6279 : _GEN_6247; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6319 = _T_1034 ? _GEN_6280 : _GEN_6248; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6320 = _T_1034 ? _GEN_6281 : _GEN_6249; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6321 = _T_1034 ? _GEN_6282 : _GEN_6250; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6322 = _T_1034 ? _GEN_6283 : _GEN_6251; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_6323 = _T_1034 ? _GEN_6284 : _GEN_6252; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [127:0] _next_reg_T_267 = $signed(_T_300) * $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:95]
  wire [63:0] _GEN_6325 = 5'h1 == rd ? _next_reg_T_267[127:64] : _GEN_6293; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6326 = 5'h2 == rd ? _next_reg_T_267[127:64] : _GEN_6294; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6327 = 5'h3 == rd ? _next_reg_T_267[127:64] : _GEN_6295; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6328 = 5'h4 == rd ? _next_reg_T_267[127:64] : _GEN_6296; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6329 = 5'h5 == rd ? _next_reg_T_267[127:64] : _GEN_6297; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6330 = 5'h6 == rd ? _next_reg_T_267[127:64] : _GEN_6298; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6331 = 5'h7 == rd ? _next_reg_T_267[127:64] : _GEN_6299; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6332 = 5'h8 == rd ? _next_reg_T_267[127:64] : _GEN_6300; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6333 = 5'h9 == rd ? _next_reg_T_267[127:64] : _GEN_6301; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6334 = 5'ha == rd ? _next_reg_T_267[127:64] : _GEN_6302; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6335 = 5'hb == rd ? _next_reg_T_267[127:64] : _GEN_6303; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6336 = 5'hc == rd ? _next_reg_T_267[127:64] : _GEN_6304; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6337 = 5'hd == rd ? _next_reg_T_267[127:64] : _GEN_6305; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6338 = 5'he == rd ? _next_reg_T_267[127:64] : _GEN_6306; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6339 = 5'hf == rd ? _next_reg_T_267[127:64] : _GEN_6307; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6340 = 5'h10 == rd ? _next_reg_T_267[127:64] : _GEN_6308; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6341 = 5'h11 == rd ? _next_reg_T_267[127:64] : _GEN_6309; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6342 = 5'h12 == rd ? _next_reg_T_267[127:64] : _GEN_6310; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6343 = 5'h13 == rd ? _next_reg_T_267[127:64] : _GEN_6311; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6344 = 5'h14 == rd ? _next_reg_T_267[127:64] : _GEN_6312; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6345 = 5'h15 == rd ? _next_reg_T_267[127:64] : _GEN_6313; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6346 = 5'h16 == rd ? _next_reg_T_267[127:64] : _GEN_6314; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6347 = 5'h17 == rd ? _next_reg_T_267[127:64] : _GEN_6315; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6348 = 5'h18 == rd ? _next_reg_T_267[127:64] : _GEN_6316; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6349 = 5'h19 == rd ? _next_reg_T_267[127:64] : _GEN_6317; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6350 = 5'h1a == rd ? _next_reg_T_267[127:64] : _GEN_6318; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6351 = 5'h1b == rd ? _next_reg_T_267[127:64] : _GEN_6319; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6352 = 5'h1c == rd ? _next_reg_T_267[127:64] : _GEN_6320; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6353 = 5'h1d == rd ? _next_reg_T_267[127:64] : _GEN_6321; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6354 = 5'h1e == rd ? _next_reg_T_267[127:64] : _GEN_6322; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6355 = 5'h1f == rd ? _next_reg_T_267[127:64] : _GEN_6323; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_6364 = _T_1041 ? _GEN_6325 : _GEN_6293; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6365 = _T_1041 ? _GEN_6326 : _GEN_6294; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6366 = _T_1041 ? _GEN_6327 : _GEN_6295; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6367 = _T_1041 ? _GEN_6328 : _GEN_6296; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6368 = _T_1041 ? _GEN_6329 : _GEN_6297; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6369 = _T_1041 ? _GEN_6330 : _GEN_6298; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6370 = _T_1041 ? _GEN_6331 : _GEN_6299; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6371 = _T_1041 ? _GEN_6332 : _GEN_6300; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6372 = _T_1041 ? _GEN_6333 : _GEN_6301; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6373 = _T_1041 ? _GEN_6334 : _GEN_6302; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6374 = _T_1041 ? _GEN_6335 : _GEN_6303; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6375 = _T_1041 ? _GEN_6336 : _GEN_6304; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6376 = _T_1041 ? _GEN_6337 : _GEN_6305; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6377 = _T_1041 ? _GEN_6338 : _GEN_6306; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6378 = _T_1041 ? _GEN_6339 : _GEN_6307; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6379 = _T_1041 ? _GEN_6340 : _GEN_6308; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6380 = _T_1041 ? _GEN_6341 : _GEN_6309; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6381 = _T_1041 ? _GEN_6342 : _GEN_6310; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6382 = _T_1041 ? _GEN_6343 : _GEN_6311; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6383 = _T_1041 ? _GEN_6344 : _GEN_6312; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6384 = _T_1041 ? _GEN_6345 : _GEN_6313; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6385 = _T_1041 ? _GEN_6346 : _GEN_6314; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6386 = _T_1041 ? _GEN_6347 : _GEN_6315; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6387 = _T_1041 ? _GEN_6348 : _GEN_6316; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6388 = _T_1041 ? _GEN_6349 : _GEN_6317; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6389 = _T_1041 ? _GEN_6350 : _GEN_6318; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6390 = _T_1041 ? _GEN_6351 : _GEN_6319; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6391 = _T_1041 ? _GEN_6352 : _GEN_6320; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6392 = _T_1041 ? _GEN_6353 : _GEN_6321; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6393 = _T_1041 ? _GEN_6354 : _GEN_6322; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_6394 = _T_1041 ? _GEN_6355 : _GEN_6323; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [64:0] _next_reg_T_270 = {1'b0,$signed(_GEN_840)}; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:72]
  wire [128:0] _next_reg_T_271 = $signed(_T_300) * $signed(_next_reg_T_270); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:72]
  wire [127:0] _next_reg_T_274 = _next_reg_T_271[127:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:88]
  wire [63:0] _GEN_6396 = 5'h1 == rd ? _next_reg_T_274[127:64] : _GEN_6364; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6397 = 5'h2 == rd ? _next_reg_T_274[127:64] : _GEN_6365; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6398 = 5'h3 == rd ? _next_reg_T_274[127:64] : _GEN_6366; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6399 = 5'h4 == rd ? _next_reg_T_274[127:64] : _GEN_6367; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6400 = 5'h5 == rd ? _next_reg_T_274[127:64] : _GEN_6368; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6401 = 5'h6 == rd ? _next_reg_T_274[127:64] : _GEN_6369; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6402 = 5'h7 == rd ? _next_reg_T_274[127:64] : _GEN_6370; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6403 = 5'h8 == rd ? _next_reg_T_274[127:64] : _GEN_6371; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6404 = 5'h9 == rd ? _next_reg_T_274[127:64] : _GEN_6372; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6405 = 5'ha == rd ? _next_reg_T_274[127:64] : _GEN_6373; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6406 = 5'hb == rd ? _next_reg_T_274[127:64] : _GEN_6374; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6407 = 5'hc == rd ? _next_reg_T_274[127:64] : _GEN_6375; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6408 = 5'hd == rd ? _next_reg_T_274[127:64] : _GEN_6376; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6409 = 5'he == rd ? _next_reg_T_274[127:64] : _GEN_6377; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6410 = 5'hf == rd ? _next_reg_T_274[127:64] : _GEN_6378; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6411 = 5'h10 == rd ? _next_reg_T_274[127:64] : _GEN_6379; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6412 = 5'h11 == rd ? _next_reg_T_274[127:64] : _GEN_6380; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6413 = 5'h12 == rd ? _next_reg_T_274[127:64] : _GEN_6381; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6414 = 5'h13 == rd ? _next_reg_T_274[127:64] : _GEN_6382; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6415 = 5'h14 == rd ? _next_reg_T_274[127:64] : _GEN_6383; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6416 = 5'h15 == rd ? _next_reg_T_274[127:64] : _GEN_6384; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6417 = 5'h16 == rd ? _next_reg_T_274[127:64] : _GEN_6385; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6418 = 5'h17 == rd ? _next_reg_T_274[127:64] : _GEN_6386; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6419 = 5'h18 == rd ? _next_reg_T_274[127:64] : _GEN_6387; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6420 = 5'h19 == rd ? _next_reg_T_274[127:64] : _GEN_6388; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6421 = 5'h1a == rd ? _next_reg_T_274[127:64] : _GEN_6389; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6422 = 5'h1b == rd ? _next_reg_T_274[127:64] : _GEN_6390; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6423 = 5'h1c == rd ? _next_reg_T_274[127:64] : _GEN_6391; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6424 = 5'h1d == rd ? _next_reg_T_274[127:64] : _GEN_6392; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6425 = 5'h1e == rd ? _next_reg_T_274[127:64] : _GEN_6393; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6426 = 5'h1f == rd ? _next_reg_T_274[127:64] : _GEN_6394; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_6435 = _T_1048 ? _GEN_6396 : _GEN_6364; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6436 = _T_1048 ? _GEN_6397 : _GEN_6365; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6437 = _T_1048 ? _GEN_6398 : _GEN_6366; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6438 = _T_1048 ? _GEN_6399 : _GEN_6367; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6439 = _T_1048 ? _GEN_6400 : _GEN_6368; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6440 = _T_1048 ? _GEN_6401 : _GEN_6369; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6441 = _T_1048 ? _GEN_6402 : _GEN_6370; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6442 = _T_1048 ? _GEN_6403 : _GEN_6371; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6443 = _T_1048 ? _GEN_6404 : _GEN_6372; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6444 = _T_1048 ? _GEN_6405 : _GEN_6373; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6445 = _T_1048 ? _GEN_6406 : _GEN_6374; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6446 = _T_1048 ? _GEN_6407 : _GEN_6375; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6447 = _T_1048 ? _GEN_6408 : _GEN_6376; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6448 = _T_1048 ? _GEN_6409 : _GEN_6377; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6449 = _T_1048 ? _GEN_6410 : _GEN_6378; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6450 = _T_1048 ? _GEN_6411 : _GEN_6379; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6451 = _T_1048 ? _GEN_6412 : _GEN_6380; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6452 = _T_1048 ? _GEN_6413 : _GEN_6381; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6453 = _T_1048 ? _GEN_6414 : _GEN_6382; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6454 = _T_1048 ? _GEN_6415 : _GEN_6383; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6455 = _T_1048 ? _GEN_6416 : _GEN_6384; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6456 = _T_1048 ? _GEN_6417 : _GEN_6385; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6457 = _T_1048 ? _GEN_6418 : _GEN_6386; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6458 = _T_1048 ? _GEN_6419 : _GEN_6387; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6459 = _T_1048 ? _GEN_6420 : _GEN_6388; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6460 = _T_1048 ? _GEN_6421 : _GEN_6389; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6461 = _T_1048 ? _GEN_6422 : _GEN_6390; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6462 = _T_1048 ? _GEN_6423 : _GEN_6391; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6463 = _T_1048 ? _GEN_6424 : _GEN_6392; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6464 = _T_1048 ? _GEN_6425 : _GEN_6393; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6465 = _T_1048 ? _GEN_6426 : _GEN_6394; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_6467 = 5'h1 == rd ? _next_reg_T_262[127:64] : _GEN_6435; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6468 = 5'h2 == rd ? _next_reg_T_262[127:64] : _GEN_6436; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6469 = 5'h3 == rd ? _next_reg_T_262[127:64] : _GEN_6437; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6470 = 5'h4 == rd ? _next_reg_T_262[127:64] : _GEN_6438; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6471 = 5'h5 == rd ? _next_reg_T_262[127:64] : _GEN_6439; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6472 = 5'h6 == rd ? _next_reg_T_262[127:64] : _GEN_6440; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6473 = 5'h7 == rd ? _next_reg_T_262[127:64] : _GEN_6441; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6474 = 5'h8 == rd ? _next_reg_T_262[127:64] : _GEN_6442; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6475 = 5'h9 == rd ? _next_reg_T_262[127:64] : _GEN_6443; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6476 = 5'ha == rd ? _next_reg_T_262[127:64] : _GEN_6444; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6477 = 5'hb == rd ? _next_reg_T_262[127:64] : _GEN_6445; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6478 = 5'hc == rd ? _next_reg_T_262[127:64] : _GEN_6446; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6479 = 5'hd == rd ? _next_reg_T_262[127:64] : _GEN_6447; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6480 = 5'he == rd ? _next_reg_T_262[127:64] : _GEN_6448; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6481 = 5'hf == rd ? _next_reg_T_262[127:64] : _GEN_6449; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6482 = 5'h10 == rd ? _next_reg_T_262[127:64] : _GEN_6450; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6483 = 5'h11 == rd ? _next_reg_T_262[127:64] : _GEN_6451; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6484 = 5'h12 == rd ? _next_reg_T_262[127:64] : _GEN_6452; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6485 = 5'h13 == rd ? _next_reg_T_262[127:64] : _GEN_6453; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6486 = 5'h14 == rd ? _next_reg_T_262[127:64] : _GEN_6454; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6487 = 5'h15 == rd ? _next_reg_T_262[127:64] : _GEN_6455; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6488 = 5'h16 == rd ? _next_reg_T_262[127:64] : _GEN_6456; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6489 = 5'h17 == rd ? _next_reg_T_262[127:64] : _GEN_6457; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6490 = 5'h18 == rd ? _next_reg_T_262[127:64] : _GEN_6458; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6491 = 5'h19 == rd ? _next_reg_T_262[127:64] : _GEN_6459; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6492 = 5'h1a == rd ? _next_reg_T_262[127:64] : _GEN_6460; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6493 = 5'h1b == rd ? _next_reg_T_262[127:64] : _GEN_6461; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6494 = 5'h1c == rd ? _next_reg_T_262[127:64] : _GEN_6462; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6495 = 5'h1d == rd ? _next_reg_T_262[127:64] : _GEN_6463; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6496 = 5'h1e == rd ? _next_reg_T_262[127:64] : _GEN_6464; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6497 = 5'h1f == rd ? _next_reg_T_262[127:64] : _GEN_6465; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_6506 = _T_1055 ? _GEN_6467 : _GEN_6435; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6507 = _T_1055 ? _GEN_6468 : _GEN_6436; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6508 = _T_1055 ? _GEN_6469 : _GEN_6437; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6509 = _T_1055 ? _GEN_6470 : _GEN_6438; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6510 = _T_1055 ? _GEN_6471 : _GEN_6439; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6511 = _T_1055 ? _GEN_6472 : _GEN_6440; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6512 = _T_1055 ? _GEN_6473 : _GEN_6441; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6513 = _T_1055 ? _GEN_6474 : _GEN_6442; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6514 = _T_1055 ? _GEN_6475 : _GEN_6443; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6515 = _T_1055 ? _GEN_6476 : _GEN_6444; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6516 = _T_1055 ? _GEN_6477 : _GEN_6445; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6517 = _T_1055 ? _GEN_6478 : _GEN_6446; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6518 = _T_1055 ? _GEN_6479 : _GEN_6447; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6519 = _T_1055 ? _GEN_6480 : _GEN_6448; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6520 = _T_1055 ? _GEN_6481 : _GEN_6449; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6521 = _T_1055 ? _GEN_6482 : _GEN_6450; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6522 = _T_1055 ? _GEN_6483 : _GEN_6451; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6523 = _T_1055 ? _GEN_6484 : _GEN_6452; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6524 = _T_1055 ? _GEN_6485 : _GEN_6453; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6525 = _T_1055 ? _GEN_6486 : _GEN_6454; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6526 = _T_1055 ? _GEN_6487 : _GEN_6455; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6527 = _T_1055 ? _GEN_6488 : _GEN_6456; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6528 = _T_1055 ? _GEN_6489 : _GEN_6457; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6529 = _T_1055 ? _GEN_6490 : _GEN_6458; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6530 = _T_1055 ? _GEN_6491 : _GEN_6459; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6531 = _T_1055 ? _GEN_6492 : _GEN_6460; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6532 = _T_1055 ? _GEN_6493 : _GEN_6461; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6533 = _T_1055 ? _GEN_6494 : _GEN_6462; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6534 = _T_1055 ? _GEN_6495 : _GEN_6463; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6535 = _T_1055 ? _GEN_6496 : _GEN_6464; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_6536 = _T_1055 ? _GEN_6497 : _GEN_6465; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [64:0] _next_reg_T_280 = $signed(_T_300) / $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 49:23]
  wire  _next_reg_T_282 = _GEN_840 == 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 51:19]
  wire [63:0] _next_reg_T_286 = 64'h0 - 64'hffffffff80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:22]
  wire  _next_reg_T_290 = _GEN_31 == _next_reg_T_286 & _GEN_840 == 64'hffffffffffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:52]
  wire [63:0] _next_reg_T_294 = _next_reg_T_290 ? _next_reg_T_286 : _next_reg_T_280[63:0]; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _next_reg_T_295 = _next_reg_T_282 ? 64'hffffffffffffffff : _next_reg_T_294; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _GEN_6538 = 5'h1 == rd ? _next_reg_T_295 : _GEN_6506; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6539 = 5'h2 == rd ? _next_reg_T_295 : _GEN_6507; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6540 = 5'h3 == rd ? _next_reg_T_295 : _GEN_6508; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6541 = 5'h4 == rd ? _next_reg_T_295 : _GEN_6509; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6542 = 5'h5 == rd ? _next_reg_T_295 : _GEN_6510; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6543 = 5'h6 == rd ? _next_reg_T_295 : _GEN_6511; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6544 = 5'h7 == rd ? _next_reg_T_295 : _GEN_6512; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6545 = 5'h8 == rd ? _next_reg_T_295 : _GEN_6513; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6546 = 5'h9 == rd ? _next_reg_T_295 : _GEN_6514; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6547 = 5'ha == rd ? _next_reg_T_295 : _GEN_6515; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6548 = 5'hb == rd ? _next_reg_T_295 : _GEN_6516; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6549 = 5'hc == rd ? _next_reg_T_295 : _GEN_6517; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6550 = 5'hd == rd ? _next_reg_T_295 : _GEN_6518; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6551 = 5'he == rd ? _next_reg_T_295 : _GEN_6519; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6552 = 5'hf == rd ? _next_reg_T_295 : _GEN_6520; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6553 = 5'h10 == rd ? _next_reg_T_295 : _GEN_6521; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6554 = 5'h11 == rd ? _next_reg_T_295 : _GEN_6522; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6555 = 5'h12 == rd ? _next_reg_T_295 : _GEN_6523; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6556 = 5'h13 == rd ? _next_reg_T_295 : _GEN_6524; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6557 = 5'h14 == rd ? _next_reg_T_295 : _GEN_6525; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6558 = 5'h15 == rd ? _next_reg_T_295 : _GEN_6526; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6559 = 5'h16 == rd ? _next_reg_T_295 : _GEN_6527; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6560 = 5'h17 == rd ? _next_reg_T_295 : _GEN_6528; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6561 = 5'h18 == rd ? _next_reg_T_295 : _GEN_6529; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6562 = 5'h19 == rd ? _next_reg_T_295 : _GEN_6530; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6563 = 5'h1a == rd ? _next_reg_T_295 : _GEN_6531; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6564 = 5'h1b == rd ? _next_reg_T_295 : _GEN_6532; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6565 = 5'h1c == rd ? _next_reg_T_295 : _GEN_6533; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6566 = 5'h1d == rd ? _next_reg_T_295 : _GEN_6534; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6567 = 5'h1e == rd ? _next_reg_T_295 : _GEN_6535; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6568 = 5'h1f == rd ? _next_reg_T_295 : _GEN_6536; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_6577 = _T_1062 ? _GEN_6538 : _GEN_6506; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6578 = _T_1062 ? _GEN_6539 : _GEN_6507; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6579 = _T_1062 ? _GEN_6540 : _GEN_6508; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6580 = _T_1062 ? _GEN_6541 : _GEN_6509; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6581 = _T_1062 ? _GEN_6542 : _GEN_6510; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6582 = _T_1062 ? _GEN_6543 : _GEN_6511; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6583 = _T_1062 ? _GEN_6544 : _GEN_6512; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6584 = _T_1062 ? _GEN_6545 : _GEN_6513; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6585 = _T_1062 ? _GEN_6546 : _GEN_6514; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6586 = _T_1062 ? _GEN_6547 : _GEN_6515; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6587 = _T_1062 ? _GEN_6548 : _GEN_6516; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6588 = _T_1062 ? _GEN_6549 : _GEN_6517; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6589 = _T_1062 ? _GEN_6550 : _GEN_6518; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6590 = _T_1062 ? _GEN_6551 : _GEN_6519; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6591 = _T_1062 ? _GEN_6552 : _GEN_6520; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6592 = _T_1062 ? _GEN_6553 : _GEN_6521; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6593 = _T_1062 ? _GEN_6554 : _GEN_6522; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6594 = _T_1062 ? _GEN_6555 : _GEN_6523; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6595 = _T_1062 ? _GEN_6556 : _GEN_6524; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6596 = _T_1062 ? _GEN_6557 : _GEN_6525; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6597 = _T_1062 ? _GEN_6558 : _GEN_6526; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6598 = _T_1062 ? _GEN_6559 : _GEN_6527; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6599 = _T_1062 ? _GEN_6560 : _GEN_6528; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6600 = _T_1062 ? _GEN_6561 : _GEN_6529; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6601 = _T_1062 ? _GEN_6562 : _GEN_6530; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6602 = _T_1062 ? _GEN_6563 : _GEN_6531; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6603 = _T_1062 ? _GEN_6564 : _GEN_6532; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6604 = _T_1062 ? _GEN_6565 : _GEN_6533; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6605 = _T_1062 ? _GEN_6566 : _GEN_6534; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6606 = _T_1062 ? _GEN_6567 : _GEN_6535; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_6607 = _T_1062 ? _GEN_6568 : _GEN_6536; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _next_reg_T_296 = _GEN_31 / _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 58:15]
  wire [63:0] _next_reg_T_299 = _next_reg_T_282 ? 64'hffffffffffffffff : _next_reg_T_296; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _GEN_6609 = 5'h1 == rd ? _next_reg_T_299 : _GEN_6577; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6610 = 5'h2 == rd ? _next_reg_T_299 : _GEN_6578; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6611 = 5'h3 == rd ? _next_reg_T_299 : _GEN_6579; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6612 = 5'h4 == rd ? _next_reg_T_299 : _GEN_6580; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6613 = 5'h5 == rd ? _next_reg_T_299 : _GEN_6581; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6614 = 5'h6 == rd ? _next_reg_T_299 : _GEN_6582; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6615 = 5'h7 == rd ? _next_reg_T_299 : _GEN_6583; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6616 = 5'h8 == rd ? _next_reg_T_299 : _GEN_6584; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6617 = 5'h9 == rd ? _next_reg_T_299 : _GEN_6585; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6618 = 5'ha == rd ? _next_reg_T_299 : _GEN_6586; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6619 = 5'hb == rd ? _next_reg_T_299 : _GEN_6587; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6620 = 5'hc == rd ? _next_reg_T_299 : _GEN_6588; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6621 = 5'hd == rd ? _next_reg_T_299 : _GEN_6589; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6622 = 5'he == rd ? _next_reg_T_299 : _GEN_6590; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6623 = 5'hf == rd ? _next_reg_T_299 : _GEN_6591; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6624 = 5'h10 == rd ? _next_reg_T_299 : _GEN_6592; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6625 = 5'h11 == rd ? _next_reg_T_299 : _GEN_6593; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6626 = 5'h12 == rd ? _next_reg_T_299 : _GEN_6594; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6627 = 5'h13 == rd ? _next_reg_T_299 : _GEN_6595; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6628 = 5'h14 == rd ? _next_reg_T_299 : _GEN_6596; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6629 = 5'h15 == rd ? _next_reg_T_299 : _GEN_6597; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6630 = 5'h16 == rd ? _next_reg_T_299 : _GEN_6598; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6631 = 5'h17 == rd ? _next_reg_T_299 : _GEN_6599; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6632 = 5'h18 == rd ? _next_reg_T_299 : _GEN_6600; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6633 = 5'h19 == rd ? _next_reg_T_299 : _GEN_6601; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6634 = 5'h1a == rd ? _next_reg_T_299 : _GEN_6602; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6635 = 5'h1b == rd ? _next_reg_T_299 : _GEN_6603; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6636 = 5'h1c == rd ? _next_reg_T_299 : _GEN_6604; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6637 = 5'h1d == rd ? _next_reg_T_299 : _GEN_6605; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6638 = 5'h1e == rd ? _next_reg_T_299 : _GEN_6606; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6639 = 5'h1f == rd ? _next_reg_T_299 : _GEN_6607; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_6648 = _T_1069 ? _GEN_6609 : _GEN_6577; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6649 = _T_1069 ? _GEN_6610 : _GEN_6578; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6650 = _T_1069 ? _GEN_6611 : _GEN_6579; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6651 = _T_1069 ? _GEN_6612 : _GEN_6580; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6652 = _T_1069 ? _GEN_6613 : _GEN_6581; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6653 = _T_1069 ? _GEN_6614 : _GEN_6582; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6654 = _T_1069 ? _GEN_6615 : _GEN_6583; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6655 = _T_1069 ? _GEN_6616 : _GEN_6584; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6656 = _T_1069 ? _GEN_6617 : _GEN_6585; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6657 = _T_1069 ? _GEN_6618 : _GEN_6586; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6658 = _T_1069 ? _GEN_6619 : _GEN_6587; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6659 = _T_1069 ? _GEN_6620 : _GEN_6588; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6660 = _T_1069 ? _GEN_6621 : _GEN_6589; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6661 = _T_1069 ? _GEN_6622 : _GEN_6590; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6662 = _T_1069 ? _GEN_6623 : _GEN_6591; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6663 = _T_1069 ? _GEN_6624 : _GEN_6592; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6664 = _T_1069 ? _GEN_6625 : _GEN_6593; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6665 = _T_1069 ? _GEN_6626 : _GEN_6594; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6666 = _T_1069 ? _GEN_6627 : _GEN_6595; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6667 = _T_1069 ? _GEN_6628 : _GEN_6596; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6668 = _T_1069 ? _GEN_6629 : _GEN_6597; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6669 = _T_1069 ? _GEN_6630 : _GEN_6598; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6670 = _T_1069 ? _GEN_6631 : _GEN_6599; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6671 = _T_1069 ? _GEN_6632 : _GEN_6600; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6672 = _T_1069 ? _GEN_6633 : _GEN_6601; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6673 = _T_1069 ? _GEN_6634 : _GEN_6602; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6674 = _T_1069 ? _GEN_6635 : _GEN_6603; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6675 = _T_1069 ? _GEN_6636 : _GEN_6604; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6676 = _T_1069 ? _GEN_6637 : _GEN_6605; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6677 = _T_1069 ? _GEN_6638 : _GEN_6606; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_6678 = _T_1069 ? _GEN_6639 : _GEN_6607; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _next_reg_T_303 = $signed(_T_300) % $signed(_T_301); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 66:42]
  wire [63:0] _next_reg_T_312 = _next_reg_T_290 ? 64'h0 : _next_reg_T_303; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _next_reg_T_313 = _next_reg_T_282 ? _GEN_31 : _next_reg_T_312; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _GEN_6680 = 5'h1 == rd ? _next_reg_T_313 : _GEN_6648; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6681 = 5'h2 == rd ? _next_reg_T_313 : _GEN_6649; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6682 = 5'h3 == rd ? _next_reg_T_313 : _GEN_6650; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6683 = 5'h4 == rd ? _next_reg_T_313 : _GEN_6651; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6684 = 5'h5 == rd ? _next_reg_T_313 : _GEN_6652; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6685 = 5'h6 == rd ? _next_reg_T_313 : _GEN_6653; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6686 = 5'h7 == rd ? _next_reg_T_313 : _GEN_6654; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6687 = 5'h8 == rd ? _next_reg_T_313 : _GEN_6655; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6688 = 5'h9 == rd ? _next_reg_T_313 : _GEN_6656; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6689 = 5'ha == rd ? _next_reg_T_313 : _GEN_6657; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6690 = 5'hb == rd ? _next_reg_T_313 : _GEN_6658; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6691 = 5'hc == rd ? _next_reg_T_313 : _GEN_6659; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6692 = 5'hd == rd ? _next_reg_T_313 : _GEN_6660; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6693 = 5'he == rd ? _next_reg_T_313 : _GEN_6661; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6694 = 5'hf == rd ? _next_reg_T_313 : _GEN_6662; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6695 = 5'h10 == rd ? _next_reg_T_313 : _GEN_6663; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6696 = 5'h11 == rd ? _next_reg_T_313 : _GEN_6664; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6697 = 5'h12 == rd ? _next_reg_T_313 : _GEN_6665; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6698 = 5'h13 == rd ? _next_reg_T_313 : _GEN_6666; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6699 = 5'h14 == rd ? _next_reg_T_313 : _GEN_6667; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6700 = 5'h15 == rd ? _next_reg_T_313 : _GEN_6668; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6701 = 5'h16 == rd ? _next_reg_T_313 : _GEN_6669; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6702 = 5'h17 == rd ? _next_reg_T_313 : _GEN_6670; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6703 = 5'h18 == rd ? _next_reg_T_313 : _GEN_6671; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6704 = 5'h19 == rd ? _next_reg_T_313 : _GEN_6672; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6705 = 5'h1a == rd ? _next_reg_T_313 : _GEN_6673; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6706 = 5'h1b == rd ? _next_reg_T_313 : _GEN_6674; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6707 = 5'h1c == rd ? _next_reg_T_313 : _GEN_6675; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6708 = 5'h1d == rd ? _next_reg_T_313 : _GEN_6676; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6709 = 5'h1e == rd ? _next_reg_T_313 : _GEN_6677; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6710 = 5'h1f == rd ? _next_reg_T_313 : _GEN_6678; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_6719 = _T_1076 ? _GEN_6680 : _GEN_6648; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6720 = _T_1076 ? _GEN_6681 : _GEN_6649; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6721 = _T_1076 ? _GEN_6682 : _GEN_6650; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6722 = _T_1076 ? _GEN_6683 : _GEN_6651; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6723 = _T_1076 ? _GEN_6684 : _GEN_6652; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6724 = _T_1076 ? _GEN_6685 : _GEN_6653; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6725 = _T_1076 ? _GEN_6686 : _GEN_6654; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6726 = _T_1076 ? _GEN_6687 : _GEN_6655; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6727 = _T_1076 ? _GEN_6688 : _GEN_6656; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6728 = _T_1076 ? _GEN_6689 : _GEN_6657; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6729 = _T_1076 ? _GEN_6690 : _GEN_6658; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6730 = _T_1076 ? _GEN_6691 : _GEN_6659; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6731 = _T_1076 ? _GEN_6692 : _GEN_6660; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6732 = _T_1076 ? _GEN_6693 : _GEN_6661; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6733 = _T_1076 ? _GEN_6694 : _GEN_6662; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6734 = _T_1076 ? _GEN_6695 : _GEN_6663; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6735 = _T_1076 ? _GEN_6696 : _GEN_6664; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6736 = _T_1076 ? _GEN_6697 : _GEN_6665; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6737 = _T_1076 ? _GEN_6698 : _GEN_6666; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6738 = _T_1076 ? _GEN_6699 : _GEN_6667; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6739 = _T_1076 ? _GEN_6700 : _GEN_6668; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6740 = _T_1076 ? _GEN_6701 : _GEN_6669; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6741 = _T_1076 ? _GEN_6702 : _GEN_6670; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6742 = _T_1076 ? _GEN_6703 : _GEN_6671; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6743 = _T_1076 ? _GEN_6704 : _GEN_6672; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6744 = _T_1076 ? _GEN_6705 : _GEN_6673; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6745 = _T_1076 ? _GEN_6706 : _GEN_6674; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6746 = _T_1076 ? _GEN_6707 : _GEN_6675; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6747 = _T_1076 ? _GEN_6708 : _GEN_6676; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6748 = _T_1076 ? _GEN_6709 : _GEN_6677; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_6749 = _T_1076 ? _GEN_6710 : _GEN_6678; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _next_reg_T_314 = _GEN_31 % _GEN_840; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 75:15]
  wire [63:0] _next_reg_T_316 = _next_reg_T_282 ? _GEN_31 : _next_reg_T_314; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _GEN_6751 = 5'h1 == rd ? _next_reg_T_316 : _GEN_6719; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6752 = 5'h2 == rd ? _next_reg_T_316 : _GEN_6720; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6753 = 5'h3 == rd ? _next_reg_T_316 : _GEN_6721; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6754 = 5'h4 == rd ? _next_reg_T_316 : _GEN_6722; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6755 = 5'h5 == rd ? _next_reg_T_316 : _GEN_6723; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6756 = 5'h6 == rd ? _next_reg_T_316 : _GEN_6724; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6757 = 5'h7 == rd ? _next_reg_T_316 : _GEN_6725; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6758 = 5'h8 == rd ? _next_reg_T_316 : _GEN_6726; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6759 = 5'h9 == rd ? _next_reg_T_316 : _GEN_6727; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6760 = 5'ha == rd ? _next_reg_T_316 : _GEN_6728; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6761 = 5'hb == rd ? _next_reg_T_316 : _GEN_6729; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6762 = 5'hc == rd ? _next_reg_T_316 : _GEN_6730; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6763 = 5'hd == rd ? _next_reg_T_316 : _GEN_6731; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6764 = 5'he == rd ? _next_reg_T_316 : _GEN_6732; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6765 = 5'hf == rd ? _next_reg_T_316 : _GEN_6733; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6766 = 5'h10 == rd ? _next_reg_T_316 : _GEN_6734; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6767 = 5'h11 == rd ? _next_reg_T_316 : _GEN_6735; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6768 = 5'h12 == rd ? _next_reg_T_316 : _GEN_6736; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6769 = 5'h13 == rd ? _next_reg_T_316 : _GEN_6737; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6770 = 5'h14 == rd ? _next_reg_T_316 : _GEN_6738; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6771 = 5'h15 == rd ? _next_reg_T_316 : _GEN_6739; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6772 = 5'h16 == rd ? _next_reg_T_316 : _GEN_6740; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6773 = 5'h17 == rd ? _next_reg_T_316 : _GEN_6741; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6774 = 5'h18 == rd ? _next_reg_T_316 : _GEN_6742; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6775 = 5'h19 == rd ? _next_reg_T_316 : _GEN_6743; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6776 = 5'h1a == rd ? _next_reg_T_316 : _GEN_6744; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6777 = 5'h1b == rd ? _next_reg_T_316 : _GEN_6745; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6778 = 5'h1c == rd ? _next_reg_T_316 : _GEN_6746; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6779 = 5'h1d == rd ? _next_reg_T_316 : _GEN_6747; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6780 = 5'h1e == rd ? _next_reg_T_316 : _GEN_6748; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6781 = 5'h1f == rd ? _next_reg_T_316 : _GEN_6749; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_6790 = _T_1083 ? _GEN_6751 : _GEN_6719; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6791 = _T_1083 ? _GEN_6752 : _GEN_6720; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6792 = _T_1083 ? _GEN_6753 : _GEN_6721; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6793 = _T_1083 ? _GEN_6754 : _GEN_6722; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6794 = _T_1083 ? _GEN_6755 : _GEN_6723; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6795 = _T_1083 ? _GEN_6756 : _GEN_6724; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6796 = _T_1083 ? _GEN_6757 : _GEN_6725; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6797 = _T_1083 ? _GEN_6758 : _GEN_6726; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6798 = _T_1083 ? _GEN_6759 : _GEN_6727; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6799 = _T_1083 ? _GEN_6760 : _GEN_6728; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6800 = _T_1083 ? _GEN_6761 : _GEN_6729; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6801 = _T_1083 ? _GEN_6762 : _GEN_6730; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6802 = _T_1083 ? _GEN_6763 : _GEN_6731; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6803 = _T_1083 ? _GEN_6764 : _GEN_6732; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6804 = _T_1083 ? _GEN_6765 : _GEN_6733; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6805 = _T_1083 ? _GEN_6766 : _GEN_6734; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6806 = _T_1083 ? _GEN_6767 : _GEN_6735; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6807 = _T_1083 ? _GEN_6768 : _GEN_6736; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6808 = _T_1083 ? _GEN_6769 : _GEN_6737; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6809 = _T_1083 ? _GEN_6770 : _GEN_6738; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6810 = _T_1083 ? _GEN_6771 : _GEN_6739; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6811 = _T_1083 ? _GEN_6772 : _GEN_6740; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6812 = _T_1083 ? _GEN_6773 : _GEN_6741; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6813 = _T_1083 ? _GEN_6774 : _GEN_6742; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6814 = _T_1083 ? _GEN_6775 : _GEN_6743; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6815 = _T_1083 ? _GEN_6776 : _GEN_6744; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6816 = _T_1083 ? _GEN_6777 : _GEN_6745; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6817 = _T_1083 ? _GEN_6778 : _GEN_6746; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6818 = _T_1083 ? _GEN_6779 : _GEN_6747; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6819 = _T_1083 ? _GEN_6780 : _GEN_6748; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_6820 = _T_1083 ? _GEN_6781 : _GEN_6749; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _next_reg_T_319 = _GEN_31[31:0] * _GEN_840[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:78]
  wire  next_reg_signBit_20 = _next_reg_T_319[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_322 = next_reg_signBit_20 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_323 = {_next_reg_T_322,_next_reg_T_319[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_6822 = 5'h1 == rd ? _next_reg_T_323 : _GEN_6790; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6823 = 5'h2 == rd ? _next_reg_T_323 : _GEN_6791; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6824 = 5'h3 == rd ? _next_reg_T_323 : _GEN_6792; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6825 = 5'h4 == rd ? _next_reg_T_323 : _GEN_6793; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6826 = 5'h5 == rd ? _next_reg_T_323 : _GEN_6794; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6827 = 5'h6 == rd ? _next_reg_T_323 : _GEN_6795; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6828 = 5'h7 == rd ? _next_reg_T_323 : _GEN_6796; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6829 = 5'h8 == rd ? _next_reg_T_323 : _GEN_6797; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6830 = 5'h9 == rd ? _next_reg_T_323 : _GEN_6798; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6831 = 5'ha == rd ? _next_reg_T_323 : _GEN_6799; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6832 = 5'hb == rd ? _next_reg_T_323 : _GEN_6800; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6833 = 5'hc == rd ? _next_reg_T_323 : _GEN_6801; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6834 = 5'hd == rd ? _next_reg_T_323 : _GEN_6802; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6835 = 5'he == rd ? _next_reg_T_323 : _GEN_6803; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6836 = 5'hf == rd ? _next_reg_T_323 : _GEN_6804; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6837 = 5'h10 == rd ? _next_reg_T_323 : _GEN_6805; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6838 = 5'h11 == rd ? _next_reg_T_323 : _GEN_6806; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6839 = 5'h12 == rd ? _next_reg_T_323 : _GEN_6807; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6840 = 5'h13 == rd ? _next_reg_T_323 : _GEN_6808; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6841 = 5'h14 == rd ? _next_reg_T_323 : _GEN_6809; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6842 = 5'h15 == rd ? _next_reg_T_323 : _GEN_6810; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6843 = 5'h16 == rd ? _next_reg_T_323 : _GEN_6811; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6844 = 5'h17 == rd ? _next_reg_T_323 : _GEN_6812; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6845 = 5'h18 == rd ? _next_reg_T_323 : _GEN_6813; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6846 = 5'h19 == rd ? _next_reg_T_323 : _GEN_6814; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6847 = 5'h1a == rd ? _next_reg_T_323 : _GEN_6815; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6848 = 5'h1b == rd ? _next_reg_T_323 : _GEN_6816; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6849 = 5'h1c == rd ? _next_reg_T_323 : _GEN_6817; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6850 = 5'h1d == rd ? _next_reg_T_323 : _GEN_6818; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6851 = 5'h1e == rd ? _next_reg_T_323 : _GEN_6819; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6852 = 5'h1f == rd ? _next_reg_T_323 : _GEN_6820; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_6861 = _T_1090 ? _GEN_6822 : _GEN_6790; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6862 = _T_1090 ? _GEN_6823 : _GEN_6791; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6863 = _T_1090 ? _GEN_6824 : _GEN_6792; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6864 = _T_1090 ? _GEN_6825 : _GEN_6793; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6865 = _T_1090 ? _GEN_6826 : _GEN_6794; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6866 = _T_1090 ? _GEN_6827 : _GEN_6795; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6867 = _T_1090 ? _GEN_6828 : _GEN_6796; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6868 = _T_1090 ? _GEN_6829 : _GEN_6797; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6869 = _T_1090 ? _GEN_6830 : _GEN_6798; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6870 = _T_1090 ? _GEN_6831 : _GEN_6799; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6871 = _T_1090 ? _GEN_6832 : _GEN_6800; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6872 = _T_1090 ? _GEN_6833 : _GEN_6801; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6873 = _T_1090 ? _GEN_6834 : _GEN_6802; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6874 = _T_1090 ? _GEN_6835 : _GEN_6803; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6875 = _T_1090 ? _GEN_6836 : _GEN_6804; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6876 = _T_1090 ? _GEN_6837 : _GEN_6805; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6877 = _T_1090 ? _GEN_6838 : _GEN_6806; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6878 = _T_1090 ? _GEN_6839 : _GEN_6807; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6879 = _T_1090 ? _GEN_6840 : _GEN_6808; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6880 = _T_1090 ? _GEN_6841 : _GEN_6809; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6881 = _T_1090 ? _GEN_6842 : _GEN_6810; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6882 = _T_1090 ? _GEN_6843 : _GEN_6811; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6883 = _T_1090 ? _GEN_6844 : _GEN_6812; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6884 = _T_1090 ? _GEN_6845 : _GEN_6813; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6885 = _T_1090 ? _GEN_6846 : _GEN_6814; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6886 = _T_1090 ? _GEN_6847 : _GEN_6815; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6887 = _T_1090 ? _GEN_6848 : _GEN_6816; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6888 = _T_1090 ? _GEN_6849 : _GEN_6817; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6889 = _T_1090 ? _GEN_6850 : _GEN_6818; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6890 = _T_1090 ? _GEN_6851 : _GEN_6819; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_6891 = _T_1090 ? _GEN_6852 : _GEN_6820; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [31:0] _next_reg_T_327 = _GEN_840[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 49:34]
  wire [32:0] _next_reg_T_328 = $signed(_next_reg_T_110) / $signed(_next_reg_T_327); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 49:23]
  wire  _next_reg_T_330 = _GEN_840[31:0] == 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 51:19]
  wire [31:0] _next_reg_T_334 = 32'h0 - 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:22]
  wire  _next_reg_T_338 = _GEN_31[31:0] == _next_reg_T_334 & _GEN_840[31:0] == 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:52]
  wire [31:0] _next_reg_T_342 = _next_reg_T_338 ? _next_reg_T_334 : _next_reg_T_328[31:0]; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _next_reg_T_343 = _next_reg_T_330 ? 32'hffffffff : _next_reg_T_342; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  next_reg_signBit_21 = _next_reg_T_343[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_345 = next_reg_signBit_21 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_346 = {_next_reg_T_345,_next_reg_T_343}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_6893 = 5'h1 == rd ? _next_reg_T_346 : _GEN_6861; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6894 = 5'h2 == rd ? _next_reg_T_346 : _GEN_6862; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6895 = 5'h3 == rd ? _next_reg_T_346 : _GEN_6863; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6896 = 5'h4 == rd ? _next_reg_T_346 : _GEN_6864; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6897 = 5'h5 == rd ? _next_reg_T_346 : _GEN_6865; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6898 = 5'h6 == rd ? _next_reg_T_346 : _GEN_6866; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6899 = 5'h7 == rd ? _next_reg_T_346 : _GEN_6867; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6900 = 5'h8 == rd ? _next_reg_T_346 : _GEN_6868; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6901 = 5'h9 == rd ? _next_reg_T_346 : _GEN_6869; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6902 = 5'ha == rd ? _next_reg_T_346 : _GEN_6870; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6903 = 5'hb == rd ? _next_reg_T_346 : _GEN_6871; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6904 = 5'hc == rd ? _next_reg_T_346 : _GEN_6872; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6905 = 5'hd == rd ? _next_reg_T_346 : _GEN_6873; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6906 = 5'he == rd ? _next_reg_T_346 : _GEN_6874; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6907 = 5'hf == rd ? _next_reg_T_346 : _GEN_6875; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6908 = 5'h10 == rd ? _next_reg_T_346 : _GEN_6876; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6909 = 5'h11 == rd ? _next_reg_T_346 : _GEN_6877; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6910 = 5'h12 == rd ? _next_reg_T_346 : _GEN_6878; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6911 = 5'h13 == rd ? _next_reg_T_346 : _GEN_6879; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6912 = 5'h14 == rd ? _next_reg_T_346 : _GEN_6880; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6913 = 5'h15 == rd ? _next_reg_T_346 : _GEN_6881; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6914 = 5'h16 == rd ? _next_reg_T_346 : _GEN_6882; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6915 = 5'h17 == rd ? _next_reg_T_346 : _GEN_6883; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6916 = 5'h18 == rd ? _next_reg_T_346 : _GEN_6884; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6917 = 5'h19 == rd ? _next_reg_T_346 : _GEN_6885; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6918 = 5'h1a == rd ? _next_reg_T_346 : _GEN_6886; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6919 = 5'h1b == rd ? _next_reg_T_346 : _GEN_6887; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6920 = 5'h1c == rd ? _next_reg_T_346 : _GEN_6888; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6921 = 5'h1d == rd ? _next_reg_T_346 : _GEN_6889; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6922 = 5'h1e == rd ? _next_reg_T_346 : _GEN_6890; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6923 = 5'h1f == rd ? _next_reg_T_346 : _GEN_6891; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_6932 = _T_1097 ? _GEN_6893 : _GEN_6861; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6933 = _T_1097 ? _GEN_6894 : _GEN_6862; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6934 = _T_1097 ? _GEN_6895 : _GEN_6863; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6935 = _T_1097 ? _GEN_6896 : _GEN_6864; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6936 = _T_1097 ? _GEN_6897 : _GEN_6865; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6937 = _T_1097 ? _GEN_6898 : _GEN_6866; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6938 = _T_1097 ? _GEN_6899 : _GEN_6867; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6939 = _T_1097 ? _GEN_6900 : _GEN_6868; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6940 = _T_1097 ? _GEN_6901 : _GEN_6869; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6941 = _T_1097 ? _GEN_6902 : _GEN_6870; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6942 = _T_1097 ? _GEN_6903 : _GEN_6871; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6943 = _T_1097 ? _GEN_6904 : _GEN_6872; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6944 = _T_1097 ? _GEN_6905 : _GEN_6873; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6945 = _T_1097 ? _GEN_6906 : _GEN_6874; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6946 = _T_1097 ? _GEN_6907 : _GEN_6875; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6947 = _T_1097 ? _GEN_6908 : _GEN_6876; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6948 = _T_1097 ? _GEN_6909 : _GEN_6877; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6949 = _T_1097 ? _GEN_6910 : _GEN_6878; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6950 = _T_1097 ? _GEN_6911 : _GEN_6879; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6951 = _T_1097 ? _GEN_6912 : _GEN_6880; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6952 = _T_1097 ? _GEN_6913 : _GEN_6881; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6953 = _T_1097 ? _GEN_6914 : _GEN_6882; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6954 = _T_1097 ? _GEN_6915 : _GEN_6883; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6955 = _T_1097 ? _GEN_6916 : _GEN_6884; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6956 = _T_1097 ? _GEN_6917 : _GEN_6885; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6957 = _T_1097 ? _GEN_6918 : _GEN_6886; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6958 = _T_1097 ? _GEN_6919 : _GEN_6887; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6959 = _T_1097 ? _GEN_6920 : _GEN_6888; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6960 = _T_1097 ? _GEN_6921 : _GEN_6889; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6961 = _T_1097 ? _GEN_6922 : _GEN_6890; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_6962 = _T_1097 ? _GEN_6923 : _GEN_6891; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [31:0] _next_reg_T_349 = _GEN_31[31:0] / _GEN_840[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 58:15]
  wire [31:0] _next_reg_T_352 = _next_reg_T_330 ? 32'hffffffff : _next_reg_T_349; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  next_reg_signBit_22 = _next_reg_T_352[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_354 = next_reg_signBit_22 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_355 = {_next_reg_T_354,_next_reg_T_352}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_6964 = 5'h1 == rd ? _next_reg_T_355 : _GEN_6932; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6965 = 5'h2 == rd ? _next_reg_T_355 : _GEN_6933; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6966 = 5'h3 == rd ? _next_reg_T_355 : _GEN_6934; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6967 = 5'h4 == rd ? _next_reg_T_355 : _GEN_6935; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6968 = 5'h5 == rd ? _next_reg_T_355 : _GEN_6936; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6969 = 5'h6 == rd ? _next_reg_T_355 : _GEN_6937; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6970 = 5'h7 == rd ? _next_reg_T_355 : _GEN_6938; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6971 = 5'h8 == rd ? _next_reg_T_355 : _GEN_6939; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6972 = 5'h9 == rd ? _next_reg_T_355 : _GEN_6940; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6973 = 5'ha == rd ? _next_reg_T_355 : _GEN_6941; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6974 = 5'hb == rd ? _next_reg_T_355 : _GEN_6942; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6975 = 5'hc == rd ? _next_reg_T_355 : _GEN_6943; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6976 = 5'hd == rd ? _next_reg_T_355 : _GEN_6944; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6977 = 5'he == rd ? _next_reg_T_355 : _GEN_6945; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6978 = 5'hf == rd ? _next_reg_T_355 : _GEN_6946; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6979 = 5'h10 == rd ? _next_reg_T_355 : _GEN_6947; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6980 = 5'h11 == rd ? _next_reg_T_355 : _GEN_6948; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6981 = 5'h12 == rd ? _next_reg_T_355 : _GEN_6949; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6982 = 5'h13 == rd ? _next_reg_T_355 : _GEN_6950; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6983 = 5'h14 == rd ? _next_reg_T_355 : _GEN_6951; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6984 = 5'h15 == rd ? _next_reg_T_355 : _GEN_6952; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6985 = 5'h16 == rd ? _next_reg_T_355 : _GEN_6953; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6986 = 5'h17 == rd ? _next_reg_T_355 : _GEN_6954; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6987 = 5'h18 == rd ? _next_reg_T_355 : _GEN_6955; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6988 = 5'h19 == rd ? _next_reg_T_355 : _GEN_6956; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6989 = 5'h1a == rd ? _next_reg_T_355 : _GEN_6957; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6990 = 5'h1b == rd ? _next_reg_T_355 : _GEN_6958; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6991 = 5'h1c == rd ? _next_reg_T_355 : _GEN_6959; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6992 = 5'h1d == rd ? _next_reg_T_355 : _GEN_6960; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6993 = 5'h1e == rd ? _next_reg_T_355 : _GEN_6961; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_6994 = 5'h1f == rd ? _next_reg_T_355 : _GEN_6962; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_7003 = _T_1104 ? _GEN_6964 : _GEN_6932; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7004 = _T_1104 ? _GEN_6965 : _GEN_6933; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7005 = _T_1104 ? _GEN_6966 : _GEN_6934; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7006 = _T_1104 ? _GEN_6967 : _GEN_6935; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7007 = _T_1104 ? _GEN_6968 : _GEN_6936; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7008 = _T_1104 ? _GEN_6969 : _GEN_6937; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7009 = _T_1104 ? _GEN_6970 : _GEN_6938; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7010 = _T_1104 ? _GEN_6971 : _GEN_6939; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7011 = _T_1104 ? _GEN_6972 : _GEN_6940; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7012 = _T_1104 ? _GEN_6973 : _GEN_6941; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7013 = _T_1104 ? _GEN_6974 : _GEN_6942; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7014 = _T_1104 ? _GEN_6975 : _GEN_6943; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7015 = _T_1104 ? _GEN_6976 : _GEN_6944; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7016 = _T_1104 ? _GEN_6977 : _GEN_6945; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7017 = _T_1104 ? _GEN_6978 : _GEN_6946; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7018 = _T_1104 ? _GEN_6979 : _GEN_6947; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7019 = _T_1104 ? _GEN_6980 : _GEN_6948; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7020 = _T_1104 ? _GEN_6981 : _GEN_6949; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7021 = _T_1104 ? _GEN_6982 : _GEN_6950; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7022 = _T_1104 ? _GEN_6983 : _GEN_6951; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7023 = _T_1104 ? _GEN_6984 : _GEN_6952; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7024 = _T_1104 ? _GEN_6985 : _GEN_6953; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7025 = _T_1104 ? _GEN_6986 : _GEN_6954; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7026 = _T_1104 ? _GEN_6987 : _GEN_6955; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7027 = _T_1104 ? _GEN_6988 : _GEN_6956; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7028 = _T_1104 ? _GEN_6989 : _GEN_6957; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7029 = _T_1104 ? _GEN_6990 : _GEN_6958; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7030 = _T_1104 ? _GEN_6991 : _GEN_6959; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7031 = _T_1104 ? _GEN_6992 : _GEN_6960; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7032 = _T_1104 ? _GEN_6993 : _GEN_6961; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_7033 = _T_1104 ? _GEN_6994 : _GEN_6962; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [31:0] _next_reg_T_361 = $signed(_next_reg_T_110) % $signed(_next_reg_T_327); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 66:42]
  wire [31:0] _next_reg_T_370 = _next_reg_T_338 ? 32'h0 : _next_reg_T_361; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _next_reg_T_371 = _next_reg_T_330 ? _GEN_31[31:0] : _next_reg_T_370; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  next_reg_signBit_23 = _next_reg_T_371[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_373 = next_reg_signBit_23 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_374 = {_next_reg_T_373,_next_reg_T_371}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_7035 = 5'h1 == rd ? _next_reg_T_374 : _GEN_7003; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7036 = 5'h2 == rd ? _next_reg_T_374 : _GEN_7004; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7037 = 5'h3 == rd ? _next_reg_T_374 : _GEN_7005; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7038 = 5'h4 == rd ? _next_reg_T_374 : _GEN_7006; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7039 = 5'h5 == rd ? _next_reg_T_374 : _GEN_7007; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7040 = 5'h6 == rd ? _next_reg_T_374 : _GEN_7008; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7041 = 5'h7 == rd ? _next_reg_T_374 : _GEN_7009; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7042 = 5'h8 == rd ? _next_reg_T_374 : _GEN_7010; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7043 = 5'h9 == rd ? _next_reg_T_374 : _GEN_7011; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7044 = 5'ha == rd ? _next_reg_T_374 : _GEN_7012; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7045 = 5'hb == rd ? _next_reg_T_374 : _GEN_7013; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7046 = 5'hc == rd ? _next_reg_T_374 : _GEN_7014; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7047 = 5'hd == rd ? _next_reg_T_374 : _GEN_7015; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7048 = 5'he == rd ? _next_reg_T_374 : _GEN_7016; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7049 = 5'hf == rd ? _next_reg_T_374 : _GEN_7017; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7050 = 5'h10 == rd ? _next_reg_T_374 : _GEN_7018; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7051 = 5'h11 == rd ? _next_reg_T_374 : _GEN_7019; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7052 = 5'h12 == rd ? _next_reg_T_374 : _GEN_7020; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7053 = 5'h13 == rd ? _next_reg_T_374 : _GEN_7021; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7054 = 5'h14 == rd ? _next_reg_T_374 : _GEN_7022; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7055 = 5'h15 == rd ? _next_reg_T_374 : _GEN_7023; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7056 = 5'h16 == rd ? _next_reg_T_374 : _GEN_7024; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7057 = 5'h17 == rd ? _next_reg_T_374 : _GEN_7025; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7058 = 5'h18 == rd ? _next_reg_T_374 : _GEN_7026; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7059 = 5'h19 == rd ? _next_reg_T_374 : _GEN_7027; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7060 = 5'h1a == rd ? _next_reg_T_374 : _GEN_7028; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7061 = 5'h1b == rd ? _next_reg_T_374 : _GEN_7029; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7062 = 5'h1c == rd ? _next_reg_T_374 : _GEN_7030; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7063 = 5'h1d == rd ? _next_reg_T_374 : _GEN_7031; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7064 = 5'h1e == rd ? _next_reg_T_374 : _GEN_7032; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7065 = 5'h1f == rd ? _next_reg_T_374 : _GEN_7033; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_7074 = _T_1111 ? _GEN_7035 : _GEN_7003; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7075 = _T_1111 ? _GEN_7036 : _GEN_7004; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7076 = _T_1111 ? _GEN_7037 : _GEN_7005; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7077 = _T_1111 ? _GEN_7038 : _GEN_7006; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7078 = _T_1111 ? _GEN_7039 : _GEN_7007; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7079 = _T_1111 ? _GEN_7040 : _GEN_7008; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7080 = _T_1111 ? _GEN_7041 : _GEN_7009; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7081 = _T_1111 ? _GEN_7042 : _GEN_7010; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7082 = _T_1111 ? _GEN_7043 : _GEN_7011; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7083 = _T_1111 ? _GEN_7044 : _GEN_7012; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7084 = _T_1111 ? _GEN_7045 : _GEN_7013; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7085 = _T_1111 ? _GEN_7046 : _GEN_7014; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7086 = _T_1111 ? _GEN_7047 : _GEN_7015; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7087 = _T_1111 ? _GEN_7048 : _GEN_7016; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7088 = _T_1111 ? _GEN_7049 : _GEN_7017; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7089 = _T_1111 ? _GEN_7050 : _GEN_7018; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7090 = _T_1111 ? _GEN_7051 : _GEN_7019; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7091 = _T_1111 ? _GEN_7052 : _GEN_7020; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7092 = _T_1111 ? _GEN_7053 : _GEN_7021; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7093 = _T_1111 ? _GEN_7054 : _GEN_7022; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7094 = _T_1111 ? _GEN_7055 : _GEN_7023; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7095 = _T_1111 ? _GEN_7056 : _GEN_7024; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7096 = _T_1111 ? _GEN_7057 : _GEN_7025; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7097 = _T_1111 ? _GEN_7058 : _GEN_7026; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7098 = _T_1111 ? _GEN_7059 : _GEN_7027; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7099 = _T_1111 ? _GEN_7060 : _GEN_7028; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7100 = _T_1111 ? _GEN_7061 : _GEN_7029; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7101 = _T_1111 ? _GEN_7062 : _GEN_7030; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7102 = _T_1111 ? _GEN_7063 : _GEN_7031; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7103 = _T_1111 ? _GEN_7064 : _GEN_7032; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_7104 = _T_1111 ? _GEN_7065 : _GEN_7033; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [31:0] _next_reg_T_377 = _GEN_31[31:0] % _GEN_840[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 75:15]
  wire [31:0] _next_reg_T_379 = _next_reg_T_330 ? _GEN_31[31:0] : _next_reg_T_377; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  next_reg_signBit_24 = _next_reg_T_379[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_381 = next_reg_signBit_24 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_382 = {_next_reg_T_381,_next_reg_T_379}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_7106 = 5'h1 == rd ? _next_reg_T_382 : _GEN_7074; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7107 = 5'h2 == rd ? _next_reg_T_382 : _GEN_7075; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7108 = 5'h3 == rd ? _next_reg_T_382 : _GEN_7076; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7109 = 5'h4 == rd ? _next_reg_T_382 : _GEN_7077; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7110 = 5'h5 == rd ? _next_reg_T_382 : _GEN_7078; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7111 = 5'h6 == rd ? _next_reg_T_382 : _GEN_7079; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7112 = 5'h7 == rd ? _next_reg_T_382 : _GEN_7080; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7113 = 5'h8 == rd ? _next_reg_T_382 : _GEN_7081; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7114 = 5'h9 == rd ? _next_reg_T_382 : _GEN_7082; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7115 = 5'ha == rd ? _next_reg_T_382 : _GEN_7083; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7116 = 5'hb == rd ? _next_reg_T_382 : _GEN_7084; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7117 = 5'hc == rd ? _next_reg_T_382 : _GEN_7085; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7118 = 5'hd == rd ? _next_reg_T_382 : _GEN_7086; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7119 = 5'he == rd ? _next_reg_T_382 : _GEN_7087; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7120 = 5'hf == rd ? _next_reg_T_382 : _GEN_7088; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7121 = 5'h10 == rd ? _next_reg_T_382 : _GEN_7089; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7122 = 5'h11 == rd ? _next_reg_T_382 : _GEN_7090; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7123 = 5'h12 == rd ? _next_reg_T_382 : _GEN_7091; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7124 = 5'h13 == rd ? _next_reg_T_382 : _GEN_7092; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7125 = 5'h14 == rd ? _next_reg_T_382 : _GEN_7093; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7126 = 5'h15 == rd ? _next_reg_T_382 : _GEN_7094; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7127 = 5'h16 == rd ? _next_reg_T_382 : _GEN_7095; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7128 = 5'h17 == rd ? _next_reg_T_382 : _GEN_7096; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7129 = 5'h18 == rd ? _next_reg_T_382 : _GEN_7097; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7130 = 5'h19 == rd ? _next_reg_T_382 : _GEN_7098; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7131 = 5'h1a == rd ? _next_reg_T_382 : _GEN_7099; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7132 = 5'h1b == rd ? _next_reg_T_382 : _GEN_7100; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7133 = 5'h1c == rd ? _next_reg_T_382 : _GEN_7101; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7134 = 5'h1d == rd ? _next_reg_T_382 : _GEN_7102; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7135 = 5'h1e == rd ? _next_reg_T_382 : _GEN_7103; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7136 = 5'h1f == rd ? _next_reg_T_382 : _GEN_7104; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_7145 = _T_1118 ? _GEN_7106 : _GEN_7074; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7146 = _T_1118 ? _GEN_7107 : _GEN_7075; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7147 = _T_1118 ? _GEN_7108 : _GEN_7076; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7148 = _T_1118 ? _GEN_7109 : _GEN_7077; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7149 = _T_1118 ? _GEN_7110 : _GEN_7078; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7150 = _T_1118 ? _GEN_7111 : _GEN_7079; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7151 = _T_1118 ? _GEN_7112 : _GEN_7080; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7152 = _T_1118 ? _GEN_7113 : _GEN_7081; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7153 = _T_1118 ? _GEN_7114 : _GEN_7082; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7154 = _T_1118 ? _GEN_7115 : _GEN_7083; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7155 = _T_1118 ? _GEN_7116 : _GEN_7084; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7156 = _T_1118 ? _GEN_7117 : _GEN_7085; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7157 = _T_1118 ? _GEN_7118 : _GEN_7086; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7158 = _T_1118 ? _GEN_7119 : _GEN_7087; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7159 = _T_1118 ? _GEN_7120 : _GEN_7088; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7160 = _T_1118 ? _GEN_7121 : _GEN_7089; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7161 = _T_1118 ? _GEN_7122 : _GEN_7090; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7162 = _T_1118 ? _GEN_7123 : _GEN_7091; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7163 = _T_1118 ? _GEN_7124 : _GEN_7092; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7164 = _T_1118 ? _GEN_7125 : _GEN_7093; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7165 = _T_1118 ? _GEN_7126 : _GEN_7094; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7166 = _T_1118 ? _GEN_7127 : _GEN_7095; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7167 = _T_1118 ? _GEN_7128 : _GEN_7096; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7168 = _T_1118 ? _GEN_7129 : _GEN_7097; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7169 = _T_1118 ? _GEN_7130 : _GEN_7098; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7170 = _T_1118 ? _GEN_7131 : _GEN_7099; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7171 = _T_1118 ? _GEN_7132 : _GEN_7100; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7172 = _T_1118 ? _GEN_7133 : _GEN_7101; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7173 = _T_1118 ? _GEN_7134 : _GEN_7102; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7174 = _T_1118 ? _GEN_7135 : _GEN_7103; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_7175 = _T_1118 ? _GEN_7136 : _GEN_7104; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire  mstatusOld_pad4 = io_now_csr_mstatus[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_sie = io_now_csr_mstatus[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_pad3 = io_now_csr_mstatus[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_mie = io_now_csr_mstatus[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_pad2 = io_now_csr_mstatus[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_spie = io_now_csr_mstatus[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_ube = io_now_csr_mstatus[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_mpie = io_now_csr_mstatus[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_spp = io_now_csr_mstatus[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] mstatusOld_vs = io_now_csr_mstatus[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] mstatusOld_mpp = io_now_csr_mstatus[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] mstatusOld_fs = io_now_csr_mstatus[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] mstatusOld_xs = io_now_csr_mstatus[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_mprv = io_now_csr_mstatus[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_sum = io_now_csr_mstatus[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_mxr = io_now_csr_mstatus[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_tvm = io_now_csr_mstatus[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_tw = io_now_csr_mstatus[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [8:0] mstatusOld_pad0 = io_now_csr_mstatus[31:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] mstatusOld_uxl = io_now_csr_mstatus[33:32]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] mstatusOld_sxl = io_now_csr_mstatus[35:34]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_sbe = io_now_csr_mstatus[36]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_mbe = io_now_csr_mstatus[37]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [24:0] mstatusOld_pad1 = io_now_csr_mstatus[62:38]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  mstatusOld_sd = io_now_csr_mstatus[63]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire [1:0] _next_internal_privilegeMode_T = {1'h0,mstatusOld_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 125:41]
  wire  mstatusNew_sie = illegalSret | illegalSModeSret ? mstatusOld_sie : mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 124:35]
  wire  mstatusNew_spie = illegalSret | illegalSModeSret ? mstatusOld_spie : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 126:35]
  wire [5:0] next_csr_mstatus_lo_lo = {mstatusNew_spie,mstatusOld_pad2,mstatusOld_mie,mstatusOld_pad3,mstatusNew_sie,
    mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  mstatusNew_spp = (illegalSret | illegalSModeSret) & mstatusOld_spp; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 127:35]
  wire [16:0] next_csr_mstatus_lo = {mstatusOld_xs,mstatusOld_fs,mstatusOld_mpp,mstatusOld_vs,mstatusNew_spp,
    mstatusOld_mpie,mstatusOld_ube,next_csr_mstatus_lo_lo}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  mstatusNew_mprv = (illegalSret | illegalSModeSret) & mstatusOld_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 128:35]
  wire [5:0] next_csr_mstatus_hi_lo = {mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,mstatusOld_mxr,mstatusOld_sum,
    mstatusNew_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [63:0] _next_csr_mstatus_T = {mstatusOld_sd,mstatusOld_pad1,mstatusOld_mbe,mstatusOld_sbe,mstatusOld_sxl,
    mstatusOld_uxl,mstatusOld_pad0,next_csr_mstatus_hi_lo,next_csr_mstatus_lo}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _GEN_7177 = illegalSret | illegalSModeSret | _GEN_3860; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_7195 = _T_1125 ? _GEN_7177 : _GEN_3860; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire  _GEN_7207 = io_now_internal_privilegeMode == 2'h3 ? _GEN_7195 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 88:48 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_7221 = _T_1132 ? _GEN_7207 : _GEN_7195; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire  _GEN_7238 = illegalInstruction | _GEN_7221; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 133:30 145:33]
  wire  raiseExceptionIntr = io_valid & _GEN_7238; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 118:36]
  wire [63:0] _delegS_T = io_now_csr_medeleg >> exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 155:24]
  wire  delegS = _delegS_T[0] & io_now_internal_privilegeMode < 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 155:39]
  wire  _T_1151 = 8'h20 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire  _T_1168 = 8'h40 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire [63:0] _GEN_7266 = 8'h40 == io_now_csr_MXLEN ? io_now_pc : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 254:35]
  wire [63:0] _GEN_7276 = 8'h20 == io_now_csr_MXLEN ? io_now_pc : _GEN_7266; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 254:35]
  wire [63:0] _GEN_7331 = delegS ? _GEN_7276 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [63:0] _GEN_7348 = raiseExceptionIntr ? _GEN_7331 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [1:0] _GEN_7179 = illegalSret | illegalSModeSret ? io_now_internal_privilegeMode : _next_internal_privilegeMode_T
    ; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 125:35]
  wire [63:0] _GEN_7183 = illegalSret | illegalSModeSret ? io_now_csr_mstatus : _next_csr_mstatus_T; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 129:35]
  wire  _GEN_7185 = illegalSret | illegalSModeSret ? _GEN_4247 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 132:25]
  wire [63:0] _GEN_7186 = illegalSret | illegalSModeSret ? _GEN_4248 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 133:25]
  wire [1:0] _GEN_7196 = _T_1125 ? _GEN_7179 : io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [63:0] _GEN_7197 = _T_1125 ? _GEN_7183 : io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire  _GEN_7199 = _T_1125 ? _GEN_7185 : _GEN_4247; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [63:0] _GEN_7200 = _T_1125 ? _GEN_7186 : _GEN_4248; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [5:0] next_csr_mstatus_lo_lo_1 = {mstatusOld_spie,mstatusOld_pad2,mstatusOld_mpie,mstatusOld_pad3,mstatusOld_sie,
    mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [16:0] next_csr_mstatus_lo_1 = {mstatusOld_xs,mstatusOld_fs,2'h3,mstatusOld_vs,mstatusOld_spp,1'h1,mstatusOld_ube
    ,next_csr_mstatus_lo_lo_1}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [5:0] next_csr_mstatus_hi_lo_1 = {mstatusOld_tsr,mstatusOld_tw,mstatusOld_tvm,mstatusOld_mxr,mstatusOld_sum,
    mstatusOld_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [63:0] _next_csr_mstatus_T_1 = {mstatusOld_sd,mstatusOld_pad1,mstatusOld_mbe,mstatusOld_sbe,mstatusOld_sxl,
    mstatusOld_uxl,mstatusOld_pad0,next_csr_mstatus_hi_lo_1,next_csr_mstatus_lo_1}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [63:0] _GEN_7306 = _T_1168 ? io_now_pc : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 186:35]
  wire [63:0] _GEN_7316 = _T_1151 ? io_now_pc : _GEN_7306; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 186:35]
  wire [63:0] _GEN_7340 = delegS ? io_now_csr_mepc : _GEN_7316; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [63:0] _GEN_7354 = raiseExceptionIntr ? _GEN_7340 : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [1:0] _GEN_7201 = io_now_internal_privilegeMode == 2'h3 ? mstatusOld_mpp : _GEN_7196; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 88:48 92:35]
  wire [63:0] _GEN_7202 = io_now_internal_privilegeMode == 2'h3 ? _next_csr_mstatus_T_1 : _GEN_7197; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:24 88:48]
  wire  _GEN_7204 = io_now_internal_privilegeMode == 2'h3 | _GEN_7199; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 103:25 88:48]
  wire [63:0] _GEN_7205 = io_now_internal_privilegeMode == 2'h3 ? io_now_csr_mepc : _GEN_7200; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 104:25 88:48]
  wire [1:0] _GEN_7215 = _T_1132 ? _GEN_7201 : _GEN_7196; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [63:0] _GEN_7216 = _T_1132 ? _GEN_7202 : _GEN_7197; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire  _GEN_7218 = _T_1132 ? _GEN_7204 : _GEN_7199; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [63:0] _GEN_7219 = _T_1132 ? _GEN_7205 : _GEN_7200; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire  _GEN_7248 = 2'h1 == io_now_csr_stvec[1:0] | _GEN_7218; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 316:29]
  wire  _GEN_7250 = 2'h0 == io_now_csr_stvec[1:0] | _GEN_7248; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 311:29]
  wire  _GEN_7273 = 8'h40 == io_now_csr_MXLEN ? _GEN_7250 : _GEN_7218; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire  _GEN_7283 = 8'h20 == io_now_csr_MXLEN ? _GEN_7250 : _GEN_7273; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire  _GEN_7291 = 2'h1 == io_now_csr_mtvec[1:0] | _GEN_7218; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 242:29]
  wire  _GEN_7293 = 2'h0 == io_now_csr_mtvec[1:0] | _GEN_7291; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 237:29]
  wire  _GEN_7313 = _T_1168 ? _GEN_7293 : _GEN_7218; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire  _GEN_7323 = _T_1151 ? _GEN_7293 : _GEN_7313; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire  _GEN_7334 = delegS ? _GEN_7283 : _GEN_7323; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire  _GEN_7351 = raiseExceptionIntr ? _GEN_7334 : _GEN_7218; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire  global_data_setpc = io_valid & _GEN_7351; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 113:21]
  wire [2:0] _next_pc_T_32 = inst[1:0] == 2'h3 ? 3'h4 : 3'h2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 154:32]
  wire [63:0] _GEN_7455 = {{61'd0}, _next_pc_T_32}; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 154:27]
  wire [63:0] _next_pc_T_34 = io_now_pc + _GEN_7455; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 154:27]
  wire [63:0] _GEN_7236 = ~global_data_setpc ? _next_pc_T_34 : _GEN_7219; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 150:30 154:17]
  wire [31:0] _next_csr_scause_T_1 = {1'h0,25'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 252:29]
  wire  mstatusNew_2_sie = delegS ? 1'h0 : mstatusOld_sie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  mstatusNew_2_spie = delegS ? mstatusOld_sie : mstatusOld_spie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  mstatusNew_2_mie = delegS & mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire [5:0] next_csr_mstatus_lo_lo_2 = {mstatusNew_2_spie,mstatusOld_pad2,mstatusNew_2_mie,mstatusOld_pad3,
    mstatusNew_2_sie,mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [1:0] _GEN_7326 = delegS ? io_now_internal_privilegeMode : {{1'd0}, mstatusOld_spp}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  mstatusNew_2_spp = _GEN_7326[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:30]
  wire  mstatusNew_2_mpie = delegS ? mstatusOld_mpie : mstatusOld_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire [1:0] mstatusNew_2_mpp = delegS ? mstatusOld_mpp : io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire [16:0] next_csr_mstatus_lo_2 = {mstatusOld_xs,mstatusOld_fs,mstatusNew_2_mpp,mstatusOld_vs,mstatusNew_2_spp,
    mstatusNew_2_mpie,mstatusOld_ube,next_csr_mstatus_lo_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [63:0] _next_csr_mstatus_T_2 = {mstatusOld_sd,mstatusOld_pad1,mstatusOld_mbe,mstatusOld_sbe,mstatusOld_sxl,
    mstatusOld_uxl,mstatusOld_pad0,next_csr_mstatus_hi_lo_1,next_csr_mstatus_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _T_1152 = 6'h2 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [31:0] _GEN_7239 = inst[1:0] != 2'h3 ? {{16'd0}, inst[15:0]} : inst; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 271:{45,62} 272:41]
  wire  _T_1155 = 6'h1 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [63:0] mem_read_addr = io_valid ? _GEN_5801 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [63:0] _GEN_7242 = 6'h4 == exceptionNO ? mem_read_addr : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29 296:26 259:35]
  wire [63:0] mem_write_addr = io_valid ? _GEN_5908 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [63:0] _GEN_7243 = 6'h6 == exceptionNO ? mem_write_addr : _GEN_7242; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29 292:26]
  wire [63:0] _GEN_7244 = 6'hb == exceptionNO ? 64'h0 : _GEN_7243; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29 288:26]
  wire [31:0] _next_pc_T_36 = {io_now_csr_stvec[31:2], 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 312:62]
  wire [31:0] _next_pc_T_38 = {26'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_7456 = {{2'd0}, io_now_csr_stvec[31:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:60]
  wire [31:0] _next_pc_T_40 = _GEN_7456 + _next_pc_T_38; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:60]
  wire [33:0] _next_pc_T_41 = {_next_pc_T_40, 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:92]
  wire [63:0] _GEN_7249 = 2'h1 == io_now_csr_stvec[1:0] ? {{30'd0}, _next_pc_T_41} : _GEN_7236; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 317:29]
  wire [63:0] _GEN_7251 = 2'h0 == io_now_csr_stvec[1:0] ? {{32'd0}, _next_pc_T_36} : _GEN_7249; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 312:29]
  wire [63:0] _next_csr_scause_T_3 = {1'h0,57'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 252:29]
  wire [63:0] _next_pc_T_43 = {io_now_csr_stvec[63:2], 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 312:62]
  wire [63:0] _next_pc_T_45 = {58'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [63:0] _GEN_7457 = {{2'd0}, io_now_csr_stvec[63:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:60]
  wire [63:0] _next_pc_T_47 = _GEN_7457 + _next_pc_T_45; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:60]
  wire [65:0] _next_pc_T_48 = {_next_pc_T_47, 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:92]
  wire [65:0] _GEN_7262 = 2'h1 == io_now_csr_stvec[1:0] ? _next_pc_T_48 : {{2'd0}, _GEN_7236}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 317:29]
  wire [65:0] _GEN_7264 = 2'h0 == io_now_csr_stvec[1:0] ? {{2'd0}, _next_pc_T_43} : _GEN_7262; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 312:29]
  wire [63:0] _GEN_7265 = 8'h40 == io_now_csr_MXLEN ? _next_csr_scause_T_3 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 252:23]
  wire [65:0] _GEN_7274 = 8'h40 == io_now_csr_MXLEN ? _GEN_7264 : {{2'd0}, _GEN_7236}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire [63:0] _GEN_7275 = 8'h20 == io_now_csr_MXLEN ? {{32'd0}, _next_csr_scause_T_1} : _GEN_7265; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 252:23]
  wire [65:0] _GEN_7284 = 8'h20 == io_now_csr_MXLEN ? {{2'd0}, _GEN_7251} : _GEN_7274; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire [63:0] _GEN_7289 = _T_1155 ? {{32'd0}, _GEN_7239} : _GEN_7244; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire [63:0] _GEN_7290 = _T_1152 ? 64'h0 : _GEN_7289; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29 199:26]
  wire [31:0] _next_pc_T_50 = {io_now_csr_mtvec[31:2], 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 238:62]
  wire [31:0] _GEN_7458 = {{2'd0}, io_now_csr_mtvec[31:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:60]
  wire [31:0] _next_pc_T_54 = _GEN_7458 + _next_pc_T_38; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:60]
  wire [33:0] _next_pc_T_55 = {_next_pc_T_54, 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:92]
  wire [63:0] _GEN_7292 = 2'h1 == io_now_csr_mtvec[1:0] ? {{30'd0}, _next_pc_T_55} : _GEN_7236; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 243:29]
  wire [63:0] _GEN_7294 = 2'h0 == io_now_csr_mtvec[1:0] ? {{32'd0}, _next_pc_T_50} : _GEN_7292; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 238:29]
  wire [63:0] _next_pc_T_57 = {io_now_csr_mtvec[63:2], 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 238:62]
  wire [63:0] _GEN_7459 = {{2'd0}, io_now_csr_mtvec[63:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:60]
  wire [63:0] _next_pc_T_61 = _GEN_7459 + _next_pc_T_45; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:60]
  wire [65:0] _next_pc_T_62 = {_next_pc_T_61, 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:92]
  wire [65:0] _GEN_7302 = 2'h1 == io_now_csr_mtvec[1:0] ? _next_pc_T_62 : {{2'd0}, _GEN_7236}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 243:29]
  wire [65:0] _GEN_7304 = 2'h0 == io_now_csr_mtvec[1:0] ? {{2'd0}, _next_pc_T_57} : _GEN_7302; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 238:29]
  wire [63:0] _GEN_7305 = _T_1168 ? _next_csr_scause_T_3 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 185:35]
  wire [63:0] _GEN_7311 = _T_1168 ? _GEN_7290 : _GEN_1925; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire [65:0] _GEN_7314 = _T_1168 ? _GEN_7304 : {{2'd0}, _GEN_7236}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire [63:0] _GEN_7315 = _T_1151 ? {{32'd0}, _next_csr_scause_T_1} : _GEN_7305; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 185:35]
  wire [63:0] _GEN_7321 = _T_1151 ? _GEN_7290 : _GEN_7311; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire [65:0] _GEN_7324 = _T_1151 ? {{2'd0}, _GEN_7294} : _GEN_7314; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire [63:0] _GEN_7330 = delegS ? _GEN_7275 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [63:0] _GEN_7347 = raiseExceptionIntr ? _GEN_7330 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [63:0] next_csr_scause = io_valid ? _GEN_7347 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [63:0] _GEN_7339 = delegS ? io_now_csr_mcause : _GEN_7315; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [63:0] _GEN_7353 = raiseExceptionIntr ? _GEN_7339 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [63:0] next_csr_mcause = io_valid ? _GEN_7353 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [63:0] _GEN_7325 = delegS ? next_csr_scause : next_csr_mcause; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 161:35 171:35]
  wire [1:0] _GEN_7329 = delegS ? 2'h1 : 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [65:0] _GEN_7335 = delegS ? _GEN_7284 : _GEN_7324; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [63:0] _GEN_7341 = delegS ? _GEN_1925 : _GEN_7321; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [63:0] _GEN_7343 = raiseExceptionIntr ? _GEN_7325 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [63:0] _GEN_7344 = raiseExceptionIntr ? io_now_pc : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30 151:25]
  wire [63:0] _GEN_7345 = raiseExceptionIntr ? {{32'd0}, inst} : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30 152:25]
  wire [1:0] _GEN_7346 = raiseExceptionIntr ? _GEN_7329 : _GEN_7215; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [63:0] _GEN_7350 = raiseExceptionIntr ? _next_csr_mstatus_T_2 : _GEN_7216; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30 181:22]
  wire [65:0] _GEN_7352 = raiseExceptionIntr ? _GEN_7335 : {{2'd0}, _GEN_7236}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [63:0] _GEN_7355 = raiseExceptionIntr ? _GEN_7341 : _GEN_1925; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [65:0] _GEN_7406 = io_valid ? _GEN_7352 : {{2'd0}, io_now_pc}; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_mem_read_valid = io_valid & _GEN_5800; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_read_addr = io_valid ? _GEN_5801 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_read_memWidth = io_valid ? _GEN_5802 : 7'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_write_valid = io_valid & _GEN_5907; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_write_addr = io_valid ? _GEN_5908 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_write_memWidth = io_valid ? _GEN_5909 : 7'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_write_data = io_valid ? _GEN_5910 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_next_reg_0 = io_valid ? 64'h0 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 148:17 111:21]
  assign io_next_reg_1 = io_valid ? _GEN_7145 : io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_2 = io_valid ? _GEN_7146 : io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_3 = io_valid ? _GEN_7147 : io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_4 = io_valid ? _GEN_7148 : io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_5 = io_valid ? _GEN_7149 : io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_6 = io_valid ? _GEN_7150 : io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_7 = io_valid ? _GEN_7151 : io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_8 = io_valid ? _GEN_7152 : io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_9 = io_valid ? _GEN_7153 : io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_10 = io_valid ? _GEN_7154 : io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_11 = io_valid ? _GEN_7155 : io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_12 = io_valid ? _GEN_7156 : io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_13 = io_valid ? _GEN_7157 : io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_14 = io_valid ? _GEN_7158 : io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_15 = io_valid ? _GEN_7159 : io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_16 = io_valid ? _GEN_7160 : io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_17 = io_valid ? _GEN_7161 : io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_18 = io_valid ? _GEN_7162 : io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_19 = io_valid ? _GEN_7163 : io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_20 = io_valid ? _GEN_7164 : io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_21 = io_valid ? _GEN_7165 : io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_22 = io_valid ? _GEN_7166 : io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_23 = io_valid ? _GEN_7167 : io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_24 = io_valid ? _GEN_7168 : io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_25 = io_valid ? _GEN_7169 : io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_26 = io_valid ? _GEN_7170 : io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_27 = io_valid ? _GEN_7171 : io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_28 = io_valid ? _GEN_7172 : io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_29 = io_valid ? _GEN_7173 : io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_30 = io_valid ? _GEN_7174 : io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_31 = io_valid ? _GEN_7175 : io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_pc = _GEN_7406[63:0]; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 18:18]
  assign io_next_csr_misa = io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mvendorid = io_now_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_marchid = io_now_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mimpid = io_now_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mhartid = io_now_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mstatus = io_valid ? _GEN_7350 : io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mscratch = io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mtvec = io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mcounteren = io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_medeleg = io_now_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mip = io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mie = io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mepc = io_valid ? _GEN_7354 : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mcause = io_valid ? _GEN_7353 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mtval = io_valid ? _GEN_7355 : io_now_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_scause = io_valid ? _GEN_7347 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_stvec = io_now_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_sepc = io_valid ? _GEN_7348 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_MXLEN = io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_internal_privilegeMode = io_valid ? _GEN_7346 : io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_event_valid = io_valid & raiseExceptionIntr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  assign io_event_cause = io_valid ? _GEN_7343 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  assign io_event_exceptionPC = io_valid ? _GEN_7344 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  assign io_event_exceptionInst = io_valid ? _GEN_7345 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
endmodule
module RiscvCore(
  input         clock,
  input         reset,
  input  [31:0] io_inst, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  input         io_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output        io_mem_read_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_mem_read_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [6:0]  io_mem_read_memWidth, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  input  [63:0] io_mem_read_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output        io_mem_write_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_mem_write_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [6:0]  io_mem_write_memWidth, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_mem_write_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_now_pc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_4, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_5, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_6, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_7, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_8, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_9, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_10, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_11, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_12, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_13, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_14, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_15, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_16, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_17, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_18, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_19, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_20, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_21, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_22, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_23, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_24, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_25, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_26, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_27, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_28, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_29, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_30, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_31, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_misa, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mvendorid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_marchid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mimpid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mhartid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mstatus, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mtvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mcounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mip, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mie, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mcause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mtval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output        io_event_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_event_cause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_event_exceptionPC, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_event_exceptionInst // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] trans_io_inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_mem_read_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_mem_read_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [6:0] trans_io_mem_read_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_mem_read_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_mem_write_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_mem_write_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [6:0] trans_io_mem_write_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_mem_write_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [1:0] trans_io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_next_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [1:0] trans_io_next_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_event_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_event_cause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_event_exceptionPC; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_event_exceptionInst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  reg [63:0] state_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [7:0] state_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [1:0] state_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  RiscvTrans trans ( // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
    .io_inst(trans_io_inst),
    .io_valid(trans_io_valid),
    .io_mem_read_valid(trans_io_mem_read_valid),
    .io_mem_read_addr(trans_io_mem_read_addr),
    .io_mem_read_memWidth(trans_io_mem_read_memWidth),
    .io_mem_read_data(trans_io_mem_read_data),
    .io_mem_write_valid(trans_io_mem_write_valid),
    .io_mem_write_addr(trans_io_mem_write_addr),
    .io_mem_write_memWidth(trans_io_mem_write_memWidth),
    .io_mem_write_data(trans_io_mem_write_data),
    .io_now_reg_0(trans_io_now_reg_0),
    .io_now_reg_1(trans_io_now_reg_1),
    .io_now_reg_2(trans_io_now_reg_2),
    .io_now_reg_3(trans_io_now_reg_3),
    .io_now_reg_4(trans_io_now_reg_4),
    .io_now_reg_5(trans_io_now_reg_5),
    .io_now_reg_6(trans_io_now_reg_6),
    .io_now_reg_7(trans_io_now_reg_7),
    .io_now_reg_8(trans_io_now_reg_8),
    .io_now_reg_9(trans_io_now_reg_9),
    .io_now_reg_10(trans_io_now_reg_10),
    .io_now_reg_11(trans_io_now_reg_11),
    .io_now_reg_12(trans_io_now_reg_12),
    .io_now_reg_13(trans_io_now_reg_13),
    .io_now_reg_14(trans_io_now_reg_14),
    .io_now_reg_15(trans_io_now_reg_15),
    .io_now_reg_16(trans_io_now_reg_16),
    .io_now_reg_17(trans_io_now_reg_17),
    .io_now_reg_18(trans_io_now_reg_18),
    .io_now_reg_19(trans_io_now_reg_19),
    .io_now_reg_20(trans_io_now_reg_20),
    .io_now_reg_21(trans_io_now_reg_21),
    .io_now_reg_22(trans_io_now_reg_22),
    .io_now_reg_23(trans_io_now_reg_23),
    .io_now_reg_24(trans_io_now_reg_24),
    .io_now_reg_25(trans_io_now_reg_25),
    .io_now_reg_26(trans_io_now_reg_26),
    .io_now_reg_27(trans_io_now_reg_27),
    .io_now_reg_28(trans_io_now_reg_28),
    .io_now_reg_29(trans_io_now_reg_29),
    .io_now_reg_30(trans_io_now_reg_30),
    .io_now_reg_31(trans_io_now_reg_31),
    .io_now_pc(trans_io_now_pc),
    .io_now_csr_misa(trans_io_now_csr_misa),
    .io_now_csr_mvendorid(trans_io_now_csr_mvendorid),
    .io_now_csr_marchid(trans_io_now_csr_marchid),
    .io_now_csr_mimpid(trans_io_now_csr_mimpid),
    .io_now_csr_mhartid(trans_io_now_csr_mhartid),
    .io_now_csr_mstatus(trans_io_now_csr_mstatus),
    .io_now_csr_mscratch(trans_io_now_csr_mscratch),
    .io_now_csr_mtvec(trans_io_now_csr_mtvec),
    .io_now_csr_mcounteren(trans_io_now_csr_mcounteren),
    .io_now_csr_medeleg(trans_io_now_csr_medeleg),
    .io_now_csr_mip(trans_io_now_csr_mip),
    .io_now_csr_mie(trans_io_now_csr_mie),
    .io_now_csr_mepc(trans_io_now_csr_mepc),
    .io_now_csr_mcause(trans_io_now_csr_mcause),
    .io_now_csr_mtval(trans_io_now_csr_mtval),
    .io_now_csr_scause(trans_io_now_csr_scause),
    .io_now_csr_stvec(trans_io_now_csr_stvec),
    .io_now_csr_sepc(trans_io_now_csr_sepc),
    .io_now_csr_MXLEN(trans_io_now_csr_MXLEN),
    .io_now_internal_privilegeMode(trans_io_now_internal_privilegeMode),
    .io_next_reg_0(trans_io_next_reg_0),
    .io_next_reg_1(trans_io_next_reg_1),
    .io_next_reg_2(trans_io_next_reg_2),
    .io_next_reg_3(trans_io_next_reg_3),
    .io_next_reg_4(trans_io_next_reg_4),
    .io_next_reg_5(trans_io_next_reg_5),
    .io_next_reg_6(trans_io_next_reg_6),
    .io_next_reg_7(trans_io_next_reg_7),
    .io_next_reg_8(trans_io_next_reg_8),
    .io_next_reg_9(trans_io_next_reg_9),
    .io_next_reg_10(trans_io_next_reg_10),
    .io_next_reg_11(trans_io_next_reg_11),
    .io_next_reg_12(trans_io_next_reg_12),
    .io_next_reg_13(trans_io_next_reg_13),
    .io_next_reg_14(trans_io_next_reg_14),
    .io_next_reg_15(trans_io_next_reg_15),
    .io_next_reg_16(trans_io_next_reg_16),
    .io_next_reg_17(trans_io_next_reg_17),
    .io_next_reg_18(trans_io_next_reg_18),
    .io_next_reg_19(trans_io_next_reg_19),
    .io_next_reg_20(trans_io_next_reg_20),
    .io_next_reg_21(trans_io_next_reg_21),
    .io_next_reg_22(trans_io_next_reg_22),
    .io_next_reg_23(trans_io_next_reg_23),
    .io_next_reg_24(trans_io_next_reg_24),
    .io_next_reg_25(trans_io_next_reg_25),
    .io_next_reg_26(trans_io_next_reg_26),
    .io_next_reg_27(trans_io_next_reg_27),
    .io_next_reg_28(trans_io_next_reg_28),
    .io_next_reg_29(trans_io_next_reg_29),
    .io_next_reg_30(trans_io_next_reg_30),
    .io_next_reg_31(trans_io_next_reg_31),
    .io_next_pc(trans_io_next_pc),
    .io_next_csr_misa(trans_io_next_csr_misa),
    .io_next_csr_mvendorid(trans_io_next_csr_mvendorid),
    .io_next_csr_marchid(trans_io_next_csr_marchid),
    .io_next_csr_mimpid(trans_io_next_csr_mimpid),
    .io_next_csr_mhartid(trans_io_next_csr_mhartid),
    .io_next_csr_mstatus(trans_io_next_csr_mstatus),
    .io_next_csr_mscratch(trans_io_next_csr_mscratch),
    .io_next_csr_mtvec(trans_io_next_csr_mtvec),
    .io_next_csr_mcounteren(trans_io_next_csr_mcounteren),
    .io_next_csr_medeleg(trans_io_next_csr_medeleg),
    .io_next_csr_mip(trans_io_next_csr_mip),
    .io_next_csr_mie(trans_io_next_csr_mie),
    .io_next_csr_mepc(trans_io_next_csr_mepc),
    .io_next_csr_mcause(trans_io_next_csr_mcause),
    .io_next_csr_mtval(trans_io_next_csr_mtval),
    .io_next_csr_scause(trans_io_next_csr_scause),
    .io_next_csr_stvec(trans_io_next_csr_stvec),
    .io_next_csr_sepc(trans_io_next_csr_sepc),
    .io_next_csr_MXLEN(trans_io_next_csr_MXLEN),
    .io_next_internal_privilegeMode(trans_io_next_internal_privilegeMode),
    .io_event_valid(trans_io_event_valid),
    .io_event_cause(trans_io_event_cause),
    .io_event_exceptionPC(trans_io_event_exceptionPC),
    .io_event_exceptionInst(trans_io_event_exceptionInst)
  );
  assign io_mem_read_valid = trans_io_mem_read_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_read_addr = trans_io_mem_read_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_read_memWidth = trans_io_mem_read_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_write_valid = trans_io_mem_write_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_write_addr = trans_io_mem_write_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_write_memWidth = trans_io_mem_write_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_write_data = trans_io_mem_write_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_now_pc = state_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_next_reg_0 = trans_io_next_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_1 = trans_io_next_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_2 = trans_io_next_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_3 = trans_io_next_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_4 = trans_io_next_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_5 = trans_io_next_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_6 = trans_io_next_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_7 = trans_io_next_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_8 = trans_io_next_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_9 = trans_io_next_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_10 = trans_io_next_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_11 = trans_io_next_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_12 = trans_io_next_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_13 = trans_io_next_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_14 = trans_io_next_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_15 = trans_io_next_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_16 = trans_io_next_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_17 = trans_io_next_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_18 = trans_io_next_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_19 = trans_io_next_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_20 = trans_io_next_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_21 = trans_io_next_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_22 = trans_io_next_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_23 = trans_io_next_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_24 = trans_io_next_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_25 = trans_io_next_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_26 = trans_io_next_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_27 = trans_io_next_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_28 = trans_io_next_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_29 = trans_io_next_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_30 = trans_io_next_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_31 = trans_io_next_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_misa = trans_io_next_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mvendorid = trans_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_marchid = trans_io_next_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mimpid = trans_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mhartid = trans_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mstatus = trans_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mscratch = trans_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mtvec = trans_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mcounteren = trans_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mip = trans_io_next_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mie = trans_io_next_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mepc = trans_io_next_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mcause = trans_io_next_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mtval = trans_io_next_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_event_valid = trans_io_event_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign io_event_cause = trans_io_event_cause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign io_event_exceptionPC = trans_io_event_exceptionPC; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign io_event_exceptionInst = trans_io_event_exceptionInst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign trans_io_inst = io_inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 192:18]
  assign trans_io_valid = io_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 193:18]
  assign trans_io_mem_read_data = io_mem_read_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign trans_io_now_reg_0 = state_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_1 = state_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_2 = state_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_3 = state_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_4 = state_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_5 = state_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_6 = state_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_7 = state_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_8 = state_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_9 = state_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_10 = state_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_11 = state_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_12 = state_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_13 = state_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_14 = state_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_15 = state_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_16 = state_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_17 = state_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_18 = state_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_19 = state_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_20 = state_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_21 = state_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_22 = state_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_23 = state_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_24 = state_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_25 = state_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_26 = state_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_27 = state_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_28 = state_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_29 = state_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_30 = state_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_31 = state_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_pc = state_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_misa = state_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mvendorid = state_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_marchid = state_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mimpid = state_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mhartid = state_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mstatus = state_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mscratch = state_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mtvec = state_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mcounteren = state_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_medeleg = state_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mip = state_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mie = state_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mepc = state_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mcause = state_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mtval = state_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_scause = state_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_stvec = state_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_sepc = state_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_MXLEN = state_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_internal_privilegeMode = state_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_0 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_0 <= trans_io_next_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_1 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_1 <= trans_io_next_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_2 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_2 <= trans_io_next_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_3 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_3 <= trans_io_next_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_4 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_4 <= trans_io_next_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_5 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_5 <= trans_io_next_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_6 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_6 <= trans_io_next_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_7 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_7 <= trans_io_next_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_8 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_8 <= trans_io_next_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_9 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_9 <= trans_io_next_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_10 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_10 <= trans_io_next_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_11 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_11 <= trans_io_next_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_12 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_12 <= trans_io_next_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_13 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_13 <= trans_io_next_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_14 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_14 <= trans_io_next_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_15 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_15 <= trans_io_next_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_16 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_16 <= trans_io_next_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_17 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_17 <= trans_io_next_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_18 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_18 <= trans_io_next_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_19 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_19 <= trans_io_next_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_20 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_20 <= trans_io_next_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_21 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_21 <= trans_io_next_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_22 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_22 <= trans_io_next_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_23 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_23 <= trans_io_next_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_24 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_24 <= trans_io_next_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_25 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_25 <= trans_io_next_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_26 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_26 <= trans_io_next_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_27 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_27 <= trans_io_next_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_28 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_28 <= trans_io_next_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_29 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_29 <= trans_io_next_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_30 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_30 <= trans_io_next_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_31 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_31 <= trans_io_next_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_pc <= 64'h80000000; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_pc <= trans_io_next_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_misa <= 64'h8000000000001104; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_misa <= trans_io_next_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mvendorid <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mvendorid <= trans_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_marchid <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_marchid <= trans_io_next_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mimpid <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mimpid <= trans_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mhartid <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mhartid <= trans_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mstatus <= 64'h1800; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mstatus <= trans_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mscratch <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mscratch <= trans_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mtvec <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mtvec <= trans_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mcounteren <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mcounteren <= trans_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_medeleg <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_medeleg <= trans_io_next_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mip <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mip <= trans_io_next_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mie <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mie <= trans_io_next_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mepc <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mepc <= trans_io_next_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mcause <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mcause <= trans_io_next_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mtval <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mtval <= trans_io_next_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_scause <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_scause <= trans_io_next_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_stvec <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_stvec <= trans_io_next_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_sepc <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_sepc <= trans_io_next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_MXLEN <= 8'h40; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_MXLEN <= trans_io_next_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_internal_privilegeMode <= 2'h3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_internal_privilegeMode <= trans_io_next_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  state_reg_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  state_reg_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  state_reg_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  state_reg_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  state_reg_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  state_reg_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  state_reg_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  state_reg_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  state_reg_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  state_reg_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  state_reg_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  state_reg_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  state_reg_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  state_reg_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  state_reg_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  state_reg_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  state_reg_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  state_reg_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  state_reg_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  state_reg_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  state_reg_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  state_reg_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  state_reg_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  state_reg_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  state_reg_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  state_reg_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  state_reg_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  state_reg_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  state_reg_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  state_reg_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  state_reg_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  state_reg_31 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  state_pc = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  state_csr_misa = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  state_csr_mvendorid = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  state_csr_marchid = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  state_csr_mimpid = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  state_csr_mhartid = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  state_csr_mstatus = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  state_csr_mscratch = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  state_csr_mtvec = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  state_csr_mcounteren = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  state_csr_medeleg = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  state_csr_mip = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  state_csr_mie = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  state_csr_mepc = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  state_csr_mcause = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  state_csr_mtval = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  state_csr_scause = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  state_csr_stvec = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  state_csr_sepc = _RAND_50[63:0];
  _RAND_51 = {1{`RANDOM}};
  state_csr_MXLEN = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  state_internal_privilegeMode = _RAND_52[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule


module CheckerWithResult(
  input         clock,
  input         reset,
  input         io_instCommit_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [31:0] io_instCommit_inst, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_instCommit_pc, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_0, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_1, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_2, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_3, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_4, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_5, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_6, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_7, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_8, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_9, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_10, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_11, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_12, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_13, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_14, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_15, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_16, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_17, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_18, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_19, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_20, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_21, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_22, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_23, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_24, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_25, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_26, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_27, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_28, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_29, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_30, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_31, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_pc, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_misa, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mvendorid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_marchid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mimpid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mhartid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mstatus, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mstatush, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mscratch, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mtvec, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mcounteren, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_medeleg, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mideleg, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mip, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mie, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mepc, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mcause, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mtval, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_cycle, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_scounteren, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_scause, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_stvec, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_sepc, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_stval, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_sscratch, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_satp, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_pmpcfg0, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_pmpcfg1, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_pmpcfg2, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_pmpcfg3, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_pmpaddr0, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_pmpaddr1, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_pmpaddr2, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_pmpaddr3, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [7:0]  io_result_csr_MXLEN, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [7:0]  io_result_csr_IALIGN, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [7:0]  io_result_csr_ILEN, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [1:0]  io_result_internal_privilegeMode, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input         io_event_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_event_intrNO, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_event_cause, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_event_exceptionPC, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_event_exceptionInst, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input         io_mem_read_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_mem_read_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [6:0]  io_mem_read_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_mem_read_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input         io_mem_write_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_mem_write_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [6:0]  io_mem_write_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_mem_write_data // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
);
  wire  specCore_clock; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire  specCore_reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [31:0] specCore_io_inst; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire  specCore_io_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire  specCore_io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_mem_read_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [6:0] specCore_io_mem_read_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_mem_read_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire  specCore_io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_mem_write_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [6:0] specCore_io_mem_write_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_mem_write_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_now_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_0; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_1; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_3; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_4; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_6; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_7; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_8; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_9; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_10; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_11; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_12; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_13; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_14; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_15; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_16; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_17; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_18; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_19; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_20; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_21; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_22; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_23; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_24; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_25; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_26; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_27; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_28; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_29; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_30; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_31; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_misa; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_marchid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mip; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mie; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mcause; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mtval; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire  specCore_io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_event_cause; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_event_exceptionPC; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_event_exceptionInst; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire  _T_2 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 102:13]
  wire  _T_4 = io_mem_read_valid | specCore_io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 103:43]
  wire  _T_17 = io_mem_write_valid | specCore_io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 108:44]
  wire  _T_218 = io_event_valid | specCore_io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 212:33]
  wire  _T_219 = io_event_valid == specCore_io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 214:32]
  wire  _GEN_1 = _T_4 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 104:15]
  wire  _GEN_8 = _T_17 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 109:15]
  wire  _GEN_17 = io_instCommit_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 198:11]
  wire  _GEN_158 = _T_218 & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 213:11]
  RiscvCore specCore ( // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
    .clock(specCore_clock),
    .reset(specCore_reset),
    .io_inst(specCore_io_inst),
    .io_valid(specCore_io_valid),
    .io_mem_read_valid(specCore_io_mem_read_valid),
    .io_mem_read_addr(specCore_io_mem_read_addr),
    .io_mem_read_memWidth(specCore_io_mem_read_memWidth),
    .io_mem_read_data(specCore_io_mem_read_data),
    .io_mem_write_valid(specCore_io_mem_write_valid),
    .io_mem_write_addr(specCore_io_mem_write_addr),
    .io_mem_write_memWidth(specCore_io_mem_write_memWidth),
    .io_mem_write_data(specCore_io_mem_write_data),
    .io_now_pc(specCore_io_now_pc),
    .io_next_reg_0(specCore_io_next_reg_0),
    .io_next_reg_1(specCore_io_next_reg_1),
    .io_next_reg_2(specCore_io_next_reg_2),
    .io_next_reg_3(specCore_io_next_reg_3),
    .io_next_reg_4(specCore_io_next_reg_4),
    .io_next_reg_5(specCore_io_next_reg_5),
    .io_next_reg_6(specCore_io_next_reg_6),
    .io_next_reg_7(specCore_io_next_reg_7),
    .io_next_reg_8(specCore_io_next_reg_8),
    .io_next_reg_9(specCore_io_next_reg_9),
    .io_next_reg_10(specCore_io_next_reg_10),
    .io_next_reg_11(specCore_io_next_reg_11),
    .io_next_reg_12(specCore_io_next_reg_12),
    .io_next_reg_13(specCore_io_next_reg_13),
    .io_next_reg_14(specCore_io_next_reg_14),
    .io_next_reg_15(specCore_io_next_reg_15),
    .io_next_reg_16(specCore_io_next_reg_16),
    .io_next_reg_17(specCore_io_next_reg_17),
    .io_next_reg_18(specCore_io_next_reg_18),
    .io_next_reg_19(specCore_io_next_reg_19),
    .io_next_reg_20(specCore_io_next_reg_20),
    .io_next_reg_21(specCore_io_next_reg_21),
    .io_next_reg_22(specCore_io_next_reg_22),
    .io_next_reg_23(specCore_io_next_reg_23),
    .io_next_reg_24(specCore_io_next_reg_24),
    .io_next_reg_25(specCore_io_next_reg_25),
    .io_next_reg_26(specCore_io_next_reg_26),
    .io_next_reg_27(specCore_io_next_reg_27),
    .io_next_reg_28(specCore_io_next_reg_28),
    .io_next_reg_29(specCore_io_next_reg_29),
    .io_next_reg_30(specCore_io_next_reg_30),
    .io_next_reg_31(specCore_io_next_reg_31),
    .io_next_csr_misa(specCore_io_next_csr_misa),
    .io_next_csr_mvendorid(specCore_io_next_csr_mvendorid),
    .io_next_csr_marchid(specCore_io_next_csr_marchid),
    .io_next_csr_mimpid(specCore_io_next_csr_mimpid),
    .io_next_csr_mhartid(specCore_io_next_csr_mhartid),
    .io_next_csr_mstatus(specCore_io_next_csr_mstatus),
    .io_next_csr_mscratch(specCore_io_next_csr_mscratch),
    .io_next_csr_mtvec(specCore_io_next_csr_mtvec),
    .io_next_csr_mcounteren(specCore_io_next_csr_mcounteren),
    .io_next_csr_mip(specCore_io_next_csr_mip),
    .io_next_csr_mie(specCore_io_next_csr_mie),
    .io_next_csr_mepc(specCore_io_next_csr_mepc),
    .io_next_csr_mcause(specCore_io_next_csr_mcause),
    .io_next_csr_mtval(specCore_io_next_csr_mtval),
    .io_event_valid(specCore_io_event_valid),
    .io_event_cause(specCore_io_event_cause),
    .io_event_exceptionPC(specCore_io_event_exceptionPC),
    .io_event_exceptionInst(specCore_io_event_exceptionInst)
  );
  assign specCore_clock = clock;
  assign specCore_reset = reset;
  assign specCore_io_inst = io_instCommit_inst; // @[src/main/scala/rvspeccore/checker/Checker.scala 89:21]
  assign specCore_io_valid = io_instCommit_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 88:21]
  assign specCore_io_mem_read_data = io_mem_read_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 113:33]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_mem_read_valid == specCore_io_mem_read_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:102 assert(regDelay(io.mem.get.read.valid) === regDelay(specCore.io.mem.read.valid))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 102:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_mem_read_valid == specCore_io_mem_read_valid)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 102:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4 & _T_2 & ~(io_mem_read_addr == specCore_io_mem_read_addr)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:104 assert(regDelay(io.mem.get.read.addr) === regDelay(specCore.io.mem.read.addr))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 104:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4 & _T_2 & ~(io_mem_read_addr == specCore_io_mem_read_addr)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 104:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1 & ~(io_mem_read_memWidth == specCore_io_mem_read_memWidth)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:105 assert(regDelay(io.mem.get.read.memWidth) === regDelay(specCore.io.mem.read.memWidth))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 105:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_1 & ~(io_mem_read_memWidth == specCore_io_mem_read_memWidth)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 105:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(io_mem_write_valid == specCore_io_mem_write_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:107 assert(regDelay(io.mem.get.write.valid) === regDelay(specCore.io.mem.write.valid))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 107:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(io_mem_write_valid == specCore_io_mem_write_valid)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 107:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_17 & _T_2 & ~(io_mem_write_addr == specCore_io_mem_write_addr)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:109 assert(regDelay(io.mem.get.write.addr) === regDelay(specCore.io.mem.write.addr))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 109:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_17 & _T_2 & ~(io_mem_write_addr == specCore_io_mem_write_addr)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 109:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_8 & ~(io_mem_write_data == specCore_io_mem_write_data)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:110 assert(regDelay(io.mem.get.write.data) === regDelay(specCore.io.mem.write.data))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 110:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_8 & ~(io_mem_write_data == specCore_io_mem_write_data)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 110:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_8 & ~(io_mem_write_memWidth == specCore_io_mem_write_memWidth)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:111 assert(regDelay(io.mem.get.write.memWidth) === regDelay(specCore.io.mem.write.memWidth))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 111:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_8 & ~(io_mem_write_memWidth == specCore_io_mem_write_memWidth)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 111:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_instCommit_valid & _T_2 & ~(io_instCommit_pc == specCore_io_now_pc)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:198 assert(regDelay(io.instCommit.pc) === regDelay(specCore.io.now.pc))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 198:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_instCommit_valid & _T_2 & ~(io_instCommit_pc == specCore_io_now_pc)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 198:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_misa == specCore_io_next_csr_misa)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_misa == specCore_io_next_csr_misa)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mvendorid == specCore_io_next_csr_mvendorid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mvendorid == specCore_io_next_csr_mvendorid)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_marchid == specCore_io_next_csr_marchid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_marchid == specCore_io_next_csr_marchid)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mimpid == specCore_io_next_csr_mimpid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mimpid == specCore_io_next_csr_mimpid)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mhartid == specCore_io_next_csr_mhartid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mhartid == specCore_io_next_csr_mhartid)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mstatus == specCore_io_next_csr_mstatus)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mstatus == specCore_io_next_csr_mstatus)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mscratch == specCore_io_next_csr_mscratch)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mscratch == specCore_io_next_csr_mscratch)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mtvec == specCore_io_next_csr_mtvec)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mtvec == specCore_io_next_csr_mtvec)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mcounteren == specCore_io_next_csr_mcounteren)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mcounteren == specCore_io_next_csr_mcounteren)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mip == specCore_io_next_csr_mip)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mip == specCore_io_next_csr_mip)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mie == specCore_io_next_csr_mie)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mie == specCore_io_next_csr_mie)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mepc == specCore_io_next_csr_mepc)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mepc == specCore_io_next_csr_mepc)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mcause == specCore_io_next_csr_mcause)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mcause == specCore_io_next_csr_mcause)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mtval == specCore_io_next_csr_mtval)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_csr_mtval == specCore_io_next_csr_mtval)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_0 == specCore_io_next_reg_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_0 == specCore_io_next_reg_0)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_1 == specCore_io_next_reg_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_1 == specCore_io_next_reg_1)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_2 == specCore_io_next_reg_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_2 == specCore_io_next_reg_2)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_3 == specCore_io_next_reg_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_3 == specCore_io_next_reg_3)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_4 == specCore_io_next_reg_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_4 == specCore_io_next_reg_4)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_5 == specCore_io_next_reg_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_5 == specCore_io_next_reg_5)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_6 == specCore_io_next_reg_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_6 == specCore_io_next_reg_6)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_7 == specCore_io_next_reg_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_7 == specCore_io_next_reg_7)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_8 == specCore_io_next_reg_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_8 == specCore_io_next_reg_8)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_9 == specCore_io_next_reg_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_9 == specCore_io_next_reg_9)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_10 == specCore_io_next_reg_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_10 == specCore_io_next_reg_10)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_11 == specCore_io_next_reg_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_11 == specCore_io_next_reg_11)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_12 == specCore_io_next_reg_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_12 == specCore_io_next_reg_12)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_13 == specCore_io_next_reg_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_13 == specCore_io_next_reg_13)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_14 == specCore_io_next_reg_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_14 == specCore_io_next_reg_14)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_15 == specCore_io_next_reg_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_15 == specCore_io_next_reg_15)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_16 == specCore_io_next_reg_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_16 == specCore_io_next_reg_16)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_17 == specCore_io_next_reg_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_17 == specCore_io_next_reg_17)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_18 == specCore_io_next_reg_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_18 == specCore_io_next_reg_18)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_19 == specCore_io_next_reg_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_19 == specCore_io_next_reg_19)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_20 == specCore_io_next_reg_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_20 == specCore_io_next_reg_20)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_21 == specCore_io_next_reg_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_21 == specCore_io_next_reg_21)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_22 == specCore_io_next_reg_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_22 == specCore_io_next_reg_22)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_23 == specCore_io_next_reg_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_23 == specCore_io_next_reg_23)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_24 == specCore_io_next_reg_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_24 == specCore_io_next_reg_24)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_25 == specCore_io_next_reg_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_25 == specCore_io_next_reg_25)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_26 == specCore_io_next_reg_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_26 == specCore_io_next_reg_26)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_27 == specCore_io_next_reg_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_27 == specCore_io_next_reg_27)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_28 == specCore_io_next_reg_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_28 == specCore_io_next_reg_28)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_29 == specCore_io_next_reg_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_29 == specCore_io_next_reg_29)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_30 == specCore_io_next_reg_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_30 == specCore_io_next_reg_30)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_31 == specCore_io_next_reg_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_17 & ~(io_result_reg_31 == specCore_io_next_reg_31)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_218 & _T_2 & ~_T_219) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Checker.scala:213 assert(\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 213:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_218 & _T_2 & ~_T_219) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 213:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_158 & ~(io_event_intrNO == 64'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:216 assert(regDelay(io.event.intrNO) === regDelay(specCore.io.event.intrNO))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 216:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_158 & ~(io_event_intrNO == 64'h0)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 216:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_158 & ~(io_event_cause == specCore_io_event_cause)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:217 assert(regDelay(io.event.cause) === regDelay(specCore.io.event.cause))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 217:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_158 & ~(io_event_cause == specCore_io_event_cause)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 217:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_158 & ~(io_event_exceptionPC == specCore_io_event_exceptionPC)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:218 assert(regDelay(io.event.exceptionPC) === regDelay(specCore.io.event.exceptionPC))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 218:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_158 & ~(io_event_exceptionPC == specCore_io_event_exceptionPC)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 218:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_158 & ~(io_event_exceptionInst == specCore_io_event_exceptionInst)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:219 assert(regDelay(io.event.exceptionInst) === regDelay(specCore.io.event.exceptionInst))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 219:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_158 & ~(io_event_exceptionInst == specCore_io_event_exceptionInst)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 219:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
