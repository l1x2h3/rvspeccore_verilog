module RiscvTrans(
  input  [31:0] io_inst, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input         io_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output        io_mem_read_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_mem_read_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [6:0]  io_mem_read_memWidth, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_mem_read_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output        io_mem_write_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_mem_write_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [6:0]  io_mem_write_memWidth, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_mem_write_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output        io_tlb_Anotherread_0_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_tlb_Anotherread_0_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_tlb_Anotherread_0_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output        io_tlb_Anotherread_1_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_tlb_Anotherread_1_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_tlb_Anotherread_1_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output        io_tlb_Anotherread_2_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_tlb_Anotherread_2_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_tlb_Anotherread_2_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_4, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_5, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_6, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_7, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_8, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_9, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_10, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_11, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_12, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_13, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_14, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_15, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_16, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_17, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_18, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_19, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_20, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_21, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_22, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_23, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_24, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_25, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_26, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_27, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_28, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_29, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_30, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_reg_31, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_pc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_misa, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mvendorid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_marchid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mimpid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mhartid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mstatus, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mtvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mcounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_medeleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mip, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mie, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mcause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_mtval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_scause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_stvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_sepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [63:0] io_now_csr_satp, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [7:0]  io_now_csr_MXLEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [7:0]  io_now_csr_IALIGN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  input  [1:0]  io_now_internal_privilegeMode, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_4, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_5, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_6, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_7, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_8, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_9, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_10, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_11, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_12, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_13, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_14, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_15, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_16, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_17, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_18, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_19, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_20, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_21, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_22, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_23, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_24, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_25, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_26, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_27, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_28, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_29, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_30, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_reg_31, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_pc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_misa, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mvendorid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_marchid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mimpid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mhartid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mstatus, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mtvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mcounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_medeleg, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mip, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mie, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mcause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_mtval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_scause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_stvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_sepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_next_csr_satp, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [7:0]  io_next_csr_MXLEN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [7:0]  io_next_csr_IALIGN, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [1:0]  io_next_internal_privilegeMode, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output        io_event_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_event_cause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_event_exceptionPC, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
  output [63:0] io_event_exceptionInst // @[src/main/scala/rvspeccore/core/RiscvCore.scala 94:14]
);
  wire  _vmEnable_T_3 = io_now_csr_satp[63:60] == 4'h8; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 110:63]
  wire  _vmEnable_T_4 = io_now_internal_privilegeMode < 2'h3; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 110:102]
  wire  vmEnable = io_now_csr_satp[63:60] == 4'h8 & io_now_internal_privilegeMode < 2'h3; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 110:71]
  wire  resultStatus = vmEnable ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 114:20 129:20]
  wire [31:0] _inst_T = resultStatus ? io_inst : 32'h13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 134:22]
  wire [31:0] inst = io_valid ? _inst_T : 32'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 134:16 112:21]
  wire [31:0] _T_1375 = inst & 32'he003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1376 = 32'h6000 == _T_1375; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  next_reg_mstatusStruct_10_mprv = io_now_csr_mstatus[17]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 60:51]
  wire [1:0] next_reg_mstatusStruct_10_mpp = io_now_csr_mstatus[12:11]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 60:51]
  wire [1:0] next_reg_pv_10 = next_reg_mstatusStruct_10_mprv ? next_reg_mstatusStruct_10_mpp :
    io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 61:30]
  wire  next_reg_vmEnable_10 = _vmEnable_T_3 & next_reg_pv_10 < 2'h3; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 62:78]
  wire [7:0] next_reg_PTE_30_flag = io_tlb_Anotherread_0_data[7:0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 275:82]
  wire  next_reg_PTEFlag_30_v = next_reg_PTE_30_flag[0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 276:42]
  wire  next_reg_PTEFlag_30_r = next_reg_PTE_30_flag[1]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 276:42]
  wire  next_reg_PTEFlag_30_w = next_reg_PTE_30_flag[2]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 276:42]
  wire  next_reg_PTEFlag_30_x = next_reg_PTE_30_flag[3]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 276:42]
  wire  _next_reg_T_758 = next_reg_PTEFlag_30_r | next_reg_PTEFlag_30_x; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 287:28]
  wire  next_reg_LevelVec_10_2_success = ~next_reg_PTEFlag_30_v | ~next_reg_PTEFlag_30_r & next_reg_PTEFlag_30_w ? 1'h0
     : _next_reg_T_758; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 277:57 284:41]
  wire  _GEN_8104 = next_reg_PTEFlag_30_r | next_reg_PTEFlag_30_x ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 287:42 291:47 299:47]
  wire  next_reg_LevelVec_10_1_valid = ~next_reg_PTEFlag_30_v | ~next_reg_PTEFlag_30_r & next_reg_PTEFlag_30_w ? 1'h0 :
    _GEN_8104; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 277:57 281:45]
  wire [7:0] next_reg_PTE_31_flag = io_tlb_Anotherread_1_data[7:0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 275:82]
  wire  next_reg_PTEFlag_31_v = next_reg_PTE_31_flag[0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 276:42]
  wire  next_reg_PTEFlag_31_r = next_reg_PTE_31_flag[1]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 276:42]
  wire  next_reg_PTEFlag_31_w = next_reg_PTE_31_flag[2]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 276:42]
  wire  next_reg_PTEFlag_31_x = next_reg_PTE_31_flag[3]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 276:42]
  wire  _next_reg_T_763 = next_reg_PTEFlag_31_r | next_reg_PTEFlag_31_x; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 287:28]
  wire  _GEN_8125 = ~next_reg_PTEFlag_31_v | ~next_reg_PTEFlag_31_r & next_reg_PTEFlag_31_w ? 1'h0 : _next_reg_T_763; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 277:57 284:41]
  wire  next_reg_LevelVec_10_1_success = next_reg_LevelVec_10_1_valid & _GEN_8125; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 271:41 319:39]
  wire  _GEN_8119 = next_reg_PTEFlag_31_r | next_reg_PTEFlag_31_x ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 287:42 291:47 299:47]
  wire  _GEN_8123 = ~next_reg_PTEFlag_31_v | ~next_reg_PTEFlag_31_r & next_reg_PTEFlag_31_w ? 1'h0 : _GEN_8119; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 277:57 281:45]
  wire  next_reg_LevelVec_10_0_valid = next_reg_LevelVec_10_1_valid & _GEN_8123; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 271:41 316:43]
  wire [7:0] next_reg_PTE_32_flag = io_tlb_Anotherread_2_data[7:0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 275:82]
  wire  next_reg_PTEFlag_32_v = next_reg_PTE_32_flag[0]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 276:42]
  wire  next_reg_PTEFlag_32_r = next_reg_PTE_32_flag[1]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 276:42]
  wire  next_reg_PTEFlag_32_w = next_reg_PTE_32_flag[2]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 276:42]
  wire  next_reg_PTEFlag_32_x = next_reg_PTE_32_flag[3]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 276:42]
  wire  _next_reg_T_768 = next_reg_PTEFlag_32_r | next_reg_PTEFlag_32_x; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 287:28]
  wire  _GEN_8136 = ~next_reg_PTEFlag_32_v | ~next_reg_PTEFlag_32_r & next_reg_PTEFlag_32_w ? 1'h0 : _next_reg_T_768; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 277:57 284:41]
  wire  next_reg_LevelVec_10_0_success = next_reg_LevelVec_10_0_valid & _GEN_8136; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 271:41 319:39]
  wire [2:0] _next_reg_successLevel_T_71 = {next_reg_LevelVec_10_2_success,next_reg_LevelVec_10_1_success,
    next_reg_LevelVec_10_0_success}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 334:39]
  wire [1:0] _next_reg_successLevel_T_73 = 3'h4 == _next_reg_successLevel_T_71 ? 2'h2 : 2'h3; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 208:25]
  wire [1:0] _next_reg_successLevel_T_75 = 3'h2 == _next_reg_successLevel_T_71 ? 2'h1 : _next_reg_successLevel_T_73; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 208:25]
  wire [1:0] next_reg_successLevel_10 = 3'h1 == _next_reg_successLevel_T_71 ? 2'h0 : _next_reg_successLevel_T_75; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 208:25]
  wire [9:0] next_reg_PTE_30_reserved = io_tlb_Anotherread_0_data[63:54]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 275:82]
  wire [43:0] next_reg_PTE_30_ppn = io_tlb_Anotherread_0_data[53:10]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 275:82]
  wire [1:0] next_reg_PTE_30_rsw = io_tlb_Anotherread_0_data[9:8]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 275:82]
  wire [63:0] _next_reg_LevelVec_2_pte_T_10 = {next_reg_PTE_30_reserved,next_reg_PTE_30_ppn,next_reg_PTE_30_rsw,
    next_reg_PTE_30_flag}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 295:50]
  wire [63:0] _GEN_8107 = next_reg_PTEFlag_30_r | next_reg_PTEFlag_30_x ? _next_reg_LevelVec_2_pte_T_10 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 287:42 295:43 309:43]
  wire [63:0] next_reg_LevelVec_10_2_pte = ~next_reg_PTEFlag_30_v | ~next_reg_PTEFlag_30_r & next_reg_PTEFlag_30_w ? 64'h0
     : _GEN_8107; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 277:57 285:41]
  wire [9:0] next_reg_PTE_31_reserved = io_tlb_Anotherread_1_data[63:54]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 275:82]
  wire [43:0] next_reg_PTE_31_ppn = io_tlb_Anotherread_1_data[53:10]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 275:82]
  wire [1:0] next_reg_PTE_31_rsw = io_tlb_Anotherread_1_data[9:8]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 275:82]
  wire [63:0] _next_reg_LevelVec_1_pte_T_10 = {next_reg_PTE_31_reserved,next_reg_PTE_31_ppn,next_reg_PTE_31_rsw,
    next_reg_PTE_31_flag}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 295:50]
  wire [63:0] _GEN_8122 = next_reg_PTEFlag_31_r | next_reg_PTEFlag_31_x ? _next_reg_LevelVec_1_pte_T_10 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 287:42 295:43 309:43]
  wire [63:0] _GEN_8126 = ~next_reg_PTEFlag_31_v | ~next_reg_PTEFlag_31_r & next_reg_PTEFlag_31_w ? 64'h0 : _GEN_8122; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 277:57 285:41]
  wire [63:0] next_reg_LevelVec_10_1_pte = next_reg_LevelVec_10_1_valid ? _GEN_8126 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 271:41 320:39]
  wire [9:0] next_reg_PTE_32_reserved = io_tlb_Anotherread_2_data[63:54]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 275:82]
  wire [43:0] next_reg_PTE_32_ppn = io_tlb_Anotherread_2_data[53:10]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 275:82]
  wire [1:0] next_reg_PTE_32_rsw = io_tlb_Anotherread_2_data[9:8]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 275:82]
  wire [63:0] _next_reg_LevelVec_0_pte_T_10 = {next_reg_PTE_32_reserved,next_reg_PTE_32_ppn,next_reg_PTE_32_rsw,
    next_reg_PTE_32_flag}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 295:50]
  wire [63:0] _GEN_8135 = next_reg_PTEFlag_32_r | next_reg_PTEFlag_32_x ? _next_reg_LevelVec_0_pte_T_10 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 287:42 295:43 309:43]
  wire [63:0] _GEN_8137 = ~next_reg_PTEFlag_32_v | ~next_reg_PTEFlag_32_r & next_reg_PTEFlag_32_w ? 64'h0 : _GEN_8135; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 277:57 285:41]
  wire [63:0] next_reg_LevelVec_10_0_pte = next_reg_LevelVec_10_0_valid ? _GEN_8137 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 271:41 320:39]
  wire [63:0] _GEN_8144 = 2'h1 == next_reg_successLevel_10 ? next_reg_LevelVec_10_1_pte : next_reg_LevelVec_10_0_pte; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 343:{48,48}]
  wire [63:0] _GEN_8145 = 2'h2 == next_reg_successLevel_10 ? next_reg_LevelVec_10_2_pte : _GEN_8144; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 343:{48,48}]
  wire  next_reg_permCheck_10 = _GEN_8145[0] & ~(next_reg_pv_10 == 2'h0 & ~_GEN_8145[4]) & ~(next_reg_pv_10 == 2'h1 &
    _GEN_8145[4] & ~io_now_csr_mstatus[18]); // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 178:58]
  wire  next_reg_mstatus_mxr_10 = io_now_csr_mstatus[19]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 174:47]
  wire  next_reg_permLoad_10 = next_reg_permCheck_10 & (_GEN_8145[1] | next_reg_mstatus_mxr_10 & _GEN_8145[3]); // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 180:31]
  wire  next_reg_permStore_10 = next_reg_permCheck_10 & _GEN_8145[2]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 181:31]
  wire [43:0] _next_reg_mask_mask_T_51 = 2'h2 == next_reg_successLevel_10 ? 44'h3ffff : 44'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 217:43]
  wire [43:0] _next_reg_mask_mask_T_53 = 2'h1 == next_reg_successLevel_10 ? 44'h1ff : _next_reg_mask_mask_T_51; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 217:43]
  wire [43:0] next_reg_mask_10 = 2'h0 == next_reg_successLevel_10 ? 44'h0 : _next_reg_mask_mask_T_53; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 217:43]
  wire [43:0] _next_reg_T_796 = next_reg_mask_10 & _GEN_8145[53:10]; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 240:11]
  wire  _next_reg_T_797 = _next_reg_T_796 != 44'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 240:18]
  wire  _GEN_8164 = _next_reg_T_797 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 349:99 351:26 360:26]
  wire  _GEN_8170 = next_reg_permLoad_10 & _GEN_8164; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 346:11 371:24]
  wire  next_reg_success_10 = ~(next_reg_successLevel_10 == 2'h3) & _GEN_8170; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 335:37 376:22]
  wire  _T_1307 = inst[11:7] != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 11:63]
  wire  _T_1308 = 32'h6002 == _T_1375 & _T_1307; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_1005 = 32'h4000 == _T_1375; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_937 = 32'h4002 == _T_1375 & _T_1307; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [31:0] _T_837 = inst & 32'h707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_838 = 32'h3003 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1786 = 32'h7073 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1743 = 32'h6073 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1709 = 32'h5073 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1667 = 32'h3073 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1625 = 32'h2073 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1592 = 32'h1073 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _T_1585 = inst & 32'hfe007fff; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1586 = 32'h12000073 == _T_1585; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1580 = 32'h10500073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1573 = 32'h30200073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1566 = 32'h10200073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _T_1558 = inst & 32'hfe00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1559 = 32'h200703b == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1552 = 32'h200603b == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1545 = 32'h200503b == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1538 = 32'h200403b == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1531 = 32'h200003b == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1524 = 32'h2007033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1517 = 32'h2006033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1510 = 32'h2005033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1503 = 32'h2004033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1496 = 32'h2003033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1489 = 32'h2002033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1482 = 32'h2001033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1475 = 32'h2000033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1452 = 32'h2001 == _T_1375 & _T_1307; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [31:0] _T_1297 = inst & 32'hef83; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1298 = 32'h1 == _T_1297; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _T_1253 = inst & 32'hf003; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_1259 = _T_1307 & inst[6:2] != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 76:105]
  wire  _T_1260 = 32'h9002 == _T_1253 & _T_1259; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_1248 = 32'h8002 == _T_1253 & _T_1259; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [5:0] _T_1195 = {inst[12],inst[6:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:14]
  wire  _T_1196 = _T_1195 != 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 17:37]
  wire  _T_1198 = _T_1307 & _T_1196; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 65:105]
  wire  _T_1199 = 32'h2 == _T_1375 & _T_1198; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_1173 = 32'h6101 == _T_1297 & _T_1196; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_1161 = 32'h1 == _T_1375 & _T_1198; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_1145 = _T_1307 & inst[11:7] != 5'h2 & _T_1196; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 44:130]
  wire  _T_1146 = 32'h6001 == _T_1375 & _T_1145; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_1128 = 32'h4001 == _T_1375 & _T_1307; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire [31:0] _T_1097 = inst & 32'hf07f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:39]
  wire  _T_1101 = 32'h9002 == _T_1097 & _T_1307; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_1092 = 32'h8002 == _T_1097 & _T_1307; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_858 = 32'h3023 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_818 = 32'h6003 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_811 = 32'h4000503b == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_804 = 32'h4000003b == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_797 = 32'h503b == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_790 = 32'h103b == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_783 = 32'h3b == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_776 = 32'h40005033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_769 = 32'h5033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_762 = 32'h1033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_756 = 32'h4000501b == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_750 = 32'h501b == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_744 = 32'h101b == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _T_737 = inst & 32'hfc00707f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_738 = 32'h40005013 == _T_737; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_732 = 32'h5013 == _T_737; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_726 = 32'h1013 == _T_737; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_720 = 32'h1b == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_714 = 32'hf == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_705 = 32'h73 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_699 = 32'h100073 == inst; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_623 = 32'h2023 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_547 = 32'h1023 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_472 = 32'h23 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_452 = 32'h5003 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_433 = 32'h4003 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_413 = 32'h2003 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_393 = 32'h1003 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_373 = 32'h3 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_346 = 32'h7063 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_317 = 32'h5063 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_290 = 32'h6063 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_261 = 32'h4063 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_234 = 32'h1063 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_207 = 32'h63 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_182 = 32'h67 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_144 = 32'h40000033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_123 = 32'h4033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_116 = 32'h6033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_109 = 32'h7033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_102 = 32'h3033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_95 = 32'h2033 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_88 = 32'h33 == _T_1558; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_56 = 32'h4013 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_50 = 32'h6013 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_44 = 32'h7013 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_38 = 32'h3013 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_32 = 32'h2013 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_26 = 32'h13 == _T_837; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [4:0] _GEN_136 = _T_26 ? inst[19:15] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 19:24]
  wire [4:0] _GEN_207 = _T_32 ? inst[19:15] : _GEN_136; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_278 = _T_38 ? inst[19:15] : _GEN_207; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_349 = _T_44 ? inst[19:15] : _GEN_278; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_420 = _T_50 ? inst[19:15] : _GEN_349; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_491 = _T_56 ? inst[19:15] : _GEN_420; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_562 = _T_726 ? inst[19:15] : _GEN_491; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_633 = _T_732 ? inst[19:15] : _GEN_562; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_704 = _T_738 ? inst[19:15] : _GEN_633; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_946 = _T_88 ? inst[19:15] : _GEN_704; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1017 = _T_95 ? inst[19:15] : _GEN_946; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1088 = _T_102 ? inst[19:15] : _GEN_1017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1159 = _T_109 ? inst[19:15] : _GEN_1088; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1230 = _T_116 ? inst[19:15] : _GEN_1159; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1301 = _T_123 ? inst[19:15] : _GEN_1230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1372 = _T_762 ? inst[19:15] : _GEN_1301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1443 = _T_769 ? inst[19:15] : _GEN_1372; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1514 = _T_144 ? inst[19:15] : _GEN_1443; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1585 = _T_776 ? inst[19:15] : _GEN_1514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1806 = _T_182 ? inst[19:15] : _GEN_1585; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1862 = _T_207 ? inst[19:15] : _GEN_1806; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1887 = _T_234 ? inst[19:15] : _GEN_1862; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1912 = _T_261 ? inst[19:15] : _GEN_1887; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1937 = _T_290 ? inst[19:15] : _GEN_1912; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1962 = _T_317 ? inst[19:15] : _GEN_1937; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1987 = _T_346 ? inst[19:15] : _GEN_1962; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2195 = _T_373 ? inst[19:15] : _GEN_1987; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2448 = _T_393 ? inst[19:15] : _GEN_2195; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2701 = _T_413 ? inst[19:15] : _GEN_2448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2905 = _T_433 ? inst[19:15] : _GEN_2701; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3158 = _T_452 ? inst[19:15] : _GEN_2905; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3331 = _T_472 ? inst[19:15] : _GEN_3158; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3491 = _T_547 ? inst[19:15] : _GEN_3331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3651 = _T_623 ? inst[19:15] : _GEN_3491; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3678 = _T_699 ? inst[19:15] : _GEN_3651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3696 = _T_705 ? inst[19:15] : _GEN_3678; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3707 = _T_714 ? inst[19:15] : _GEN_3696; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3746 = _T_720 ? inst[19:15] : _GEN_3707; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3817 = _T_726 ? inst[19:15] : _GEN_3746; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3888 = _T_732 ? inst[19:15] : _GEN_3817; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3959 = _T_738 ? inst[19:15] : _GEN_3888; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4030 = _T_744 ? inst[19:15] : _GEN_3959; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4101 = _T_750 ? inst[19:15] : _GEN_4030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4172 = _T_756 ? inst[19:15] : _GEN_4101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4244 = _T_762 ? inst[19:15] : _GEN_4172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4315 = _T_769 ? inst[19:15] : _GEN_4244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4386 = _T_776 ? inst[19:15] : _GEN_4315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4457 = _T_783 ? inst[19:15] : _GEN_4386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4528 = _T_790 ? inst[19:15] : _GEN_4457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4599 = _T_797 ? inst[19:15] : _GEN_4528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4670 = _T_804 ? inst[19:15] : _GEN_4599; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4741 = _T_811 ? inst[19:15] : _GEN_4670; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4974 = _T_818 ? inst[19:15] : _GEN_4741; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5227 = _T_838 ? inst[19:15] : _GEN_4974; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5418 = _T_858 ? inst[19:15] : _GEN_5227; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5590 = _T_937 ? inst[11:7] : _GEN_5418; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6236 = _T_1092 ? inst[11:7] : _GEN_5590; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6244 = _T_1101 ? inst[11:7] : _GEN_6236; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6374 = _T_1128 ? inst[11:7] : _GEN_6244; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6446 = _T_1146 ? inst[11:7] : _GEN_6374; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6549 = _T_1161 ? inst[11:7] : _GEN_6446; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6588 = _T_1173 ? inst[11:7] : _GEN_6549; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 220:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6697 = _T_1199 ? inst[11:7] : _GEN_6588; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7080 = _T_1248 ? inst[11:7] : _GEN_6697; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7150 = _T_1260 ? inst[11:7] : _GEN_7080; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7729 = _T_1298 ? inst[11:7] : _GEN_7150; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 259:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7880 = _T_1308 ? inst[11:7] : _GEN_7729; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_8544 = _T_1452 ? inst[11:7] : _GEN_7880; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_8886 = _T_1475 ? inst[19:15] : _GEN_8544; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_8957 = _T_1482 ? inst[19:15] : _GEN_8886; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9028 = _T_1489 ? inst[19:15] : _GEN_8957; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9099 = _T_1496 ? inst[19:15] : _GEN_9028; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9170 = _T_1503 ? inst[19:15] : _GEN_9099; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9241 = _T_1510 ? inst[19:15] : _GEN_9170; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9312 = _T_1517 ? inst[19:15] : _GEN_9241; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9383 = _T_1524 ? inst[19:15] : _GEN_9312; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9454 = _T_1531 ? inst[19:15] : _GEN_9383; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9525 = _T_1538 ? inst[19:15] : _GEN_9454; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9596 = _T_1545 ? inst[19:15] : _GEN_9525; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9667 = _T_1552 ? inst[19:15] : _GEN_9596; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9738 = _T_1559 ? inst[19:15] : _GEN_9667; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9787 = _T_1566 ? inst[19:15] : _GEN_9738; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9808 = _T_1573 ? inst[19:15] : _GEN_9787; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9822 = _T_1580 ? inst[19:15] : _GEN_9808; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9829 = _T_1586 ? inst[19:15] : _GEN_9822; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9976 = _T_1592 ? inst[19:15] : _GEN_9829; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_10156 = _T_1625 ? inst[19:15] : _GEN_9976; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_10336 = _T_1667 ? inst[19:15] : _GEN_10156; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_10528 = _T_1709 ? inst[19:15] : _GEN_10336; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_10708 = _T_1743 ? inst[19:15] : _GEN_10528; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_10888 = _T_1786 ? inst[19:15] : _GEN_10708; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] rs1 = io_valid ? _GEN_10888 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 19:24]
  wire [63:0] _GEN_71 = 5'h1 == rs1 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_72 = 5'h2 == rs1 ? io_now_reg_2 : _GEN_71; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_73 = 5'h3 == rs1 ? io_now_reg_3 : _GEN_72; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_74 = 5'h4 == rs1 ? io_now_reg_4 : _GEN_73; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_75 = 5'h5 == rs1 ? io_now_reg_5 : _GEN_74; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_76 = 5'h6 == rs1 ? io_now_reg_6 : _GEN_75; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_77 = 5'h7 == rs1 ? io_now_reg_7 : _GEN_76; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_78 = 5'h8 == rs1 ? io_now_reg_8 : _GEN_77; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_79 = 5'h9 == rs1 ? io_now_reg_9 : _GEN_78; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_80 = 5'ha == rs1 ? io_now_reg_10 : _GEN_79; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_81 = 5'hb == rs1 ? io_now_reg_11 : _GEN_80; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_82 = 5'hc == rs1 ? io_now_reg_12 : _GEN_81; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_83 = 5'hd == rs1 ? io_now_reg_13 : _GEN_82; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_84 = 5'he == rs1 ? io_now_reg_14 : _GEN_83; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_85 = 5'hf == rs1 ? io_now_reg_15 : _GEN_84; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_86 = 5'h10 == rs1 ? io_now_reg_16 : _GEN_85; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_87 = 5'h11 == rs1 ? io_now_reg_17 : _GEN_86; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_88 = 5'h12 == rs1 ? io_now_reg_18 : _GEN_87; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_89 = 5'h13 == rs1 ? io_now_reg_19 : _GEN_88; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_90 = 5'h14 == rs1 ? io_now_reg_20 : _GEN_89; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_91 = 5'h15 == rs1 ? io_now_reg_21 : _GEN_90; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_92 = 5'h16 == rs1 ? io_now_reg_22 : _GEN_91; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_93 = 5'h17 == rs1 ? io_now_reg_23 : _GEN_92; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_94 = 5'h18 == rs1 ? io_now_reg_24 : _GEN_93; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_95 = 5'h19 == rs1 ? io_now_reg_25 : _GEN_94; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_96 = 5'h1a == rs1 ? io_now_reg_26 : _GEN_95; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_97 = 5'h1b == rs1 ? io_now_reg_27 : _GEN_96; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_98 = 5'h1c == rs1 ? io_now_reg_28 : _GEN_97; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_99 = 5'h1d == rs1 ? io_now_reg_29 : _GEN_98; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_100 = 5'h1e == rs1 ? io_now_reg_30 : _GEN_99; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [63:0] _GEN_101 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{63,63}]
  wire [11:0] _GEN_135 = _T_26 ? inst[31:20] : 12'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 38:27]
  wire [11:0] _GEN_206 = _T_32 ? inst[31:20] : _GEN_135; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_277 = _T_38 ? inst[31:20] : _GEN_206; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_348 = _T_44 ? inst[31:20] : _GEN_277; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_419 = _T_50 ? inst[31:20] : _GEN_348; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_490 = _T_56 ? inst[31:20] : _GEN_419; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_561 = _T_726 ? inst[31:20] : _GEN_490; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_632 = _T_732 ? inst[31:20] : _GEN_561; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_703 = _T_738 ? inst[31:20] : _GEN_632; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_1805 = _T_182 ? inst[31:20] : _GEN_703; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2194 = _T_373 ? inst[31:20] : _GEN_1805; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2447 = _T_393 ? inst[31:20] : _GEN_2194; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2700 = _T_413 ? inst[31:20] : _GEN_2447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_2904 = _T_433 ? inst[31:20] : _GEN_2700; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_3157 = _T_452 ? inst[31:20] : _GEN_2904; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_3677 = _T_699 ? inst[31:20] : _GEN_3157; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_3695 = _T_705 ? inst[31:20] : _GEN_3677; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_3706 = _T_714 ? inst[31:20] : _GEN_3695; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_3745 = _T_720 ? inst[31:20] : _GEN_3706; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_3816 = _T_726 ? inst[31:20] : _GEN_3745; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_3887 = _T_732 ? inst[31:20] : _GEN_3816; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_3958 = _T_738 ? inst[31:20] : _GEN_3887; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_4029 = _T_744 ? inst[31:20] : _GEN_3958; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_4100 = _T_750 ? inst[31:20] : _GEN_4029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_4171 = _T_756 ? inst[31:20] : _GEN_4100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_4973 = _T_818 ? inst[31:20] : _GEN_4171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_5226 = _T_838 ? inst[31:20] : _GEN_4973; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_9786 = _T_1566 ? inst[31:20] : _GEN_5226; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_9807 = _T_1573 ? inst[31:20] : _GEN_9786; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_9821 = _T_1580 ? inst[31:20] : _GEN_9807; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_9828 = _T_1586 ? inst[31:20] : _GEN_9821; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_9975 = _T_1592 ? inst[31:20] : _GEN_9828; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_10155 = _T_1625 ? inst[31:20] : _GEN_9975; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_10335 = _T_1667 ? inst[31:20] : _GEN_10155; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_10527 = _T_1709 ? inst[31:20] : _GEN_10335; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_10707 = _T_1743 ? inst[31:20] : _GEN_10527; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] _GEN_10887 = _T_1786 ? inst[31:20] : _GEN_10707; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [11:0] imm_11_0 = io_valid ? _GEN_10887 : 12'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 38:27]
  wire  imm_signBit_56 = imm_11_0[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [51:0] _imm_T_338 = imm_signBit_56 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _imm_T_339 = {_imm_T_338,imm_11_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [5:0] _imm_T_306 = {inst[12],inst[6],inst[5],inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 83:10]
  wire  imm_signBit_46 = _imm_T_306[5]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [57:0] _imm_T_308 = imm_signBit_46 ? 58'h3ffffffffffffff : 58'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _imm_T_309 = {_imm_T_308,inst[12],inst[6],inst[5],inst[4],inst[3],inst[2]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  _T_1385 = 32'he000 == _T_1375; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [63:0] _imm_T_299 = {56'h0,inst[6],inst[5],inst[12],inst[11],inst[10],3'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire  _T_1315 = 32'he002 == _T_1375; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [63:0] _imm_T_283 = {55'h0,inst[9],inst[8],inst[7],inst[12],inst[11],inst[10],3'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [63:0] _imm_T_274 = {55'h0,inst[4],inst[3],inst[2],inst[12],inst[6],inst[5],3'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _T_1233 = inst & 32'hec03; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1234 = 32'h8801 == _T_1233; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1226 = 32'h8401 == _T_1233 & _T_1196; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_1212 = 32'h8001 == _T_1233 & _T_1196; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _T_1116 = 32'he001 == _T_1375; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [8:0] _imm_T_221 = {inst[12],inst[6],inst[5],inst[2],inst[11],inst[10],inst[4],inst[3],1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire  imm_signBit_43 = _imm_T_221[8]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [54:0] _imm_T_223 = imm_signBit_43 ? 55'h7fffffffffffff : 55'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _imm_T_224 = {_imm_T_223,inst[12],inst[6],inst[5],inst[2],inst[11],inst[10],inst[4],inst[3],1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  _T_1107 = 32'hc001 == _T_1375; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [4:0] imm_lo_12 = {inst[2],inst[11],inst[5],inst[4],inst[3]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:14]
  wire [11:0] _imm_T_195 = {inst[12],inst[8],inst[10],inst[9],inst[6],inst[7],imm_lo_12,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire  imm_signBit_41 = _imm_T_195[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [51:0] _imm_T_197 = imm_signBit_41 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _imm_T_198 = {_imm_T_197,inst[12],inst[8],inst[10],inst[9],inst[6],inst[7],imm_lo_12,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  _T_1078 = 32'ha001 == _T_1375; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1014 = 32'hc000 == _T_1375; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [63:0] _imm_T_166 = {57'h0,inst[5],inst[12],inst[11],inst[10],inst[6],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire  _T_944 = 32'hc002 == _T_1375; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [63:0] _imm_T_150 = {56'h0,inst[8],inst[7],inst[12],inst[11],inst[10],inst[9],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [63:0] _imm_T_141 = {56'h0,inst[3],inst[2],inst[12],inst[6],inst[5],inst[4],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [6:0] _GEN_3329 = _T_472 ? inst[31:25] : 7'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:27]
  wire [6:0] _GEN_3489 = _T_547 ? inst[31:25] : _GEN_3329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_3649 = _T_623 ? inst[31:25] : _GEN_3489; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] _GEN_5416 = _T_858 ? inst[31:25] : _GEN_3649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [6:0] imm_11_5 = io_valid ? _GEN_5416 : 7'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:27]
  wire [4:0] _GEN_3333 = _T_472 ? inst[11:7] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:62]
  wire [4:0] _GEN_3493 = _T_547 ? inst[11:7] : _GEN_3333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3653 = _T_623 ? inst[11:7] : _GEN_3493; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5420 = _T_858 ? inst[11:7] : _GEN_3653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] imm_4_0 = io_valid ? _GEN_5420 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 39:62]
  wire [11:0] _imm_T_129 = {imm_11_5,imm_4_0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:141]
  wire  imm_signBit_39 = _imm_T_129[11]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [51:0] _imm_T_131 = imm_signBit_39 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _imm_T_132 = {_imm_T_131,imm_11_5,imm_4_0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  _GEN_1859 = _T_207 & inst[31]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:27]
  wire  _GEN_1884 = _T_234 ? inst[31] : _GEN_1859; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1909 = _T_261 ? inst[31] : _GEN_1884; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1934 = _T_290 ? inst[31] : _GEN_1909; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1959 = _T_317 ? inst[31] : _GEN_1934; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1984 = _T_346 ? inst[31] : _GEN_1959; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  imm_12 = io_valid & _GEN_1984; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:27]
  wire [31:0] _T_157 = inst & 32'h7f; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_158 = 32'h6f == _T_157; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _GEN_1693 = _T_158 & inst[20]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:132]
  wire  _GEN_1865 = _T_207 ? inst[7] : _GEN_1693; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1890 = _T_234 ? inst[7] : _GEN_1865; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1915 = _T_261 ? inst[7] : _GEN_1890; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1940 = _T_290 ? inst[7] : _GEN_1915; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1965 = _T_317 ? inst[7] : _GEN_1940; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  _GEN_1990 = _T_346 ? inst[7] : _GEN_1965; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire  imm_11 = io_valid & _GEN_1990; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:132]
  wire [5:0] _GEN_1860 = _T_207 ? inst[30:25] : 6'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:62]
  wire [5:0] _GEN_1885 = _T_234 ? inst[30:25] : _GEN_1860; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_1910 = _T_261 ? inst[30:25] : _GEN_1885; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_1935 = _T_290 ? inst[30:25] : _GEN_1910; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_1960 = _T_317 ? inst[30:25] : _GEN_1935; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] _GEN_1985 = _T_346 ? inst[30:25] : _GEN_1960; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [5:0] imm_10_5 = io_valid ? _GEN_1985 : 6'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:62]
  wire [3:0] _GEN_1864 = _T_207 ? inst[11:8] : 4'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:99]
  wire [3:0] _GEN_1889 = _T_234 ? inst[11:8] : _GEN_1864; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] _GEN_1914 = _T_261 ? inst[11:8] : _GEN_1889; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] _GEN_1939 = _T_290 ? inst[11:8] : _GEN_1914; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] _GEN_1964 = _T_317 ? inst[11:8] : _GEN_1939; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] _GEN_1989 = _T_346 ? inst[11:8] : _GEN_1964; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [3:0] imm_4_1 = io_valid ? _GEN_1989 : 4'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 40:99]
  wire [12:0] _imm_T_62 = {imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:141]
  wire  imm_signBit_18 = _imm_T_62[12]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [50:0] _imm_T_64 = imm_signBit_18 ? 51'h7ffffffffffff : 51'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _imm_T_65 = {_imm_T_64,imm_12,imm_11,imm_10_5,imm_4_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  _GEN_1691 = _T_158 & inst[31]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:27]
  wire  imm_20 = io_valid & _GEN_1691; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:27]
  wire [7:0] _GEN_1694 = _T_158 ? inst[19:12] : 8'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:99]
  wire [7:0] imm_19_12 = io_valid ? _GEN_1694 : 8'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:99]
  wire [9:0] _GEN_1692 = _T_158 ? inst[30:21] : 10'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:62]
  wire [9:0] imm_10_1 = io_valid ? _GEN_1692 : 10'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 42:62]
  wire [20:0] _imm_T_35 = {imm_20,imm_19_12,imm_11,imm_10_1,1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 52:141]
  wire  imm_signBit_11 = _imm_T_35[20]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [42:0] _imm_T_37 = imm_signBit_11 ? 43'h7ffffffffff : 43'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _imm_T_38 = {_imm_T_37,imm_20,imm_19_12,imm_11,imm_10_1,1'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire  _T_84 = 32'h17 == _T_157; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_80 = 32'h37 == _T_157; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [19:0] _GEN_774 = _T_80 ? inst[31:12] : 20'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 41:27]
  wire [19:0] _GEN_843 = _T_84 ? inst[31:12] : _GEN_774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [19:0] imm_31_12 = io_valid ? _GEN_843 : 20'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 41:27]
  wire [31:0] _imm_T_31 = {imm_31_12,12'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:141]
  wire  imm_signBit_10 = _imm_T_31[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _imm_T_33 = imm_signBit_10 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _imm_T_34 = {_imm_T_33,imm_31_12,12'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_140 = _T_26 ? _imm_T_339 : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 22:24]
  wire [63:0] _GEN_211 = _T_32 ? _imm_T_339 : _GEN_140; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_282 = _T_38 ? _imm_T_339 : _GEN_211; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_353 = _T_44 ? _imm_T_339 : _GEN_282; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_424 = _T_50 ? _imm_T_339 : _GEN_353; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_495 = _T_56 ? _imm_T_339 : _GEN_424; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_566 = _T_726 ? _imm_T_339 : _GEN_495; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_637 = _T_732 ? _imm_T_339 : _GEN_566; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_708 = _T_738 ? _imm_T_339 : _GEN_637; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_777 = _T_80 ? _imm_T_34 : _GEN_708; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:127]
  wire [63:0] _GEN_846 = _T_84 ? _imm_T_34 : _GEN_777; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 51:127]
  wire [63:0] _GEN_1697 = _T_158 ? _imm_T_38 : _GEN_846; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 52:127]
  wire [63:0] _GEN_1810 = _T_182 ? _imm_T_339 : _GEN_1697; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_1867 = _T_207 ? _imm_T_65 : _GEN_1810; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [63:0] _GEN_1892 = _T_234 ? _imm_T_65 : _GEN_1867; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [63:0] _GEN_1917 = _T_261 ? _imm_T_65 : _GEN_1892; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [63:0] _GEN_1942 = _T_290 ? _imm_T_65 : _GEN_1917; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [63:0] _GEN_1967 = _T_317 ? _imm_T_65 : _GEN_1942; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [63:0] _GEN_1992 = _T_346 ? _imm_T_65 : _GEN_1967; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 50:127]
  wire [63:0] _GEN_2199 = _T_373 ? _imm_T_339 : _GEN_1992; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_2452 = _T_393 ? _imm_T_339 : _GEN_2199; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_2705 = _T_413 ? _imm_T_339 : _GEN_2452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_2909 = _T_433 ? _imm_T_339 : _GEN_2705; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_3162 = _T_452 ? _imm_T_339 : _GEN_2909; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_3335 = _T_472 ? _imm_T_132 : _GEN_3162; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:127]
  wire [63:0] _GEN_3495 = _T_547 ? _imm_T_132 : _GEN_3335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:127]
  wire [63:0] _GEN_3655 = _T_623 ? _imm_T_132 : _GEN_3495; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:127]
  wire [63:0] _GEN_3682 = _T_699 ? _imm_T_339 : _GEN_3655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_3700 = _T_705 ? _imm_T_339 : _GEN_3682; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_3711 = _T_714 ? _imm_T_339 : _GEN_3700; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_3750 = _T_720 ? _imm_T_339 : _GEN_3711; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_3821 = _T_726 ? _imm_T_339 : _GEN_3750; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_3892 = _T_732 ? _imm_T_339 : _GEN_3821; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_3963 = _T_738 ? _imm_T_339 : _GEN_3892; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_4034 = _T_744 ? _imm_T_339 : _GEN_3963; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_4105 = _T_750 ? _imm_T_339 : _GEN_4034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_4176 = _T_756 ? _imm_T_339 : _GEN_4105; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_4978 = _T_818 ? _imm_T_339 : _GEN_4176; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_5231 = _T_838 ? _imm_T_339 : _GEN_4978; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_5422 = _T_858 ? _imm_T_132 : _GEN_5231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 49:127]
  wire [63:0] _GEN_5594 = _T_937 ? _imm_T_141 : _GEN_5422; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 140:20]
  wire [63:0] _GEN_5762 = _T_944 ? _imm_T_150 : _GEN_5594; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 145:11]
  wire [63:0] _GEN_5965 = _T_1005 ? _imm_T_166 : _GEN_5762; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 151:28]
  wire [63:0] _GEN_6199 = _T_1014 ? _imm_T_166 : _GEN_5965; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 156:11]
  wire [63:0] _GEN_6223 = _T_1078 ? _imm_T_198 : _GEN_6199; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 160:21 162:25]
  wire [63:0] _GEN_6292 = _T_1107 ? _imm_T_224 : _GEN_6223; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24 188:11]
  wire [63:0] _GEN_6336 = _T_1116 ? _imm_T_224 : _GEN_6292; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24 196:11]
  wire [63:0] _GEN_6378 = _T_1128 ? _imm_T_309 : _GEN_6336; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22 206:20]
  wire [63:0] _GEN_6701 = _T_1199 ? {{58'd0}, _imm_T_306} : _GEN_6378; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24 232:20]
  wire [63:0] _GEN_6805 = _T_1212 ? {{58'd0}, _imm_T_306} : _GEN_6701; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24 237:28]
  wire [63:0] _GEN_6909 = _T_1226 ? {{58'd0}, _imm_T_306} : _GEN_6805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24 242:28]
  wire [63:0] _GEN_7013 = _T_1234 ? _imm_T_309 : _GEN_6909; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24 247:28]
  wire [63:0] _GEN_7884 = _T_1308 ? _imm_T_274 : _GEN_7013; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24 269:20]
  wire [63:0] _GEN_8052 = _T_1315 ? _imm_T_283 : _GEN_7884; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24 274:11]
  wire [63:0] _GEN_8255 = _T_1376 ? _imm_T_299 : _GEN_8052; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22 280:28]
  wire [63:0] _GEN_8489 = _T_1385 ? _imm_T_299 : _GEN_8255; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22 285:11]
  wire [63:0] _GEN_8548 = _T_1452 ? _imm_T_309 : _GEN_8489; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25 292:20]
  wire [63:0] _GEN_9791 = _T_1566 ? _imm_T_339 : _GEN_8548; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [63:0] _GEN_9812 = _T_1573 ? _imm_T_339 : _GEN_9791; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [63:0] _GEN_9826 = _T_1580 ? _imm_T_339 : _GEN_9812; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28]
  wire [63:0] _GEN_9833 = _T_1586 ? _imm_T_339 : _GEN_9826; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28]
  wire [63:0] _GEN_9980 = _T_1592 ? _imm_T_339 : _GEN_9833; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10160 = _T_1625 ? _imm_T_339 : _GEN_9980; // @[src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10340 = _T_1667 ? _imm_T_339 : _GEN_10160; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_10532 = _T_1709 ? _imm_T_339 : _GEN_10340; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_10712 = _T_1743 ? _imm_T_339 : _GEN_10532; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] _GEN_10892 = _T_1786 ? _imm_T_339 : _GEN_10712; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 48:127]
  wire [63:0] imm = io_valid ? _GEN_10892 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 22:24]
  wire [63:0] _T_844 = _GEN_101 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:47]
  wire  _T_850 = _T_844[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_848 = _T_844[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_846 = ~_T_844[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _GEN_2092 = next_reg_success_10 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30 144:33]
  wire  _GEN_2108 = next_reg_vmEnable_10 & _GEN_2092; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_2215 = _T_373 & _GEN_2108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_2345 = next_reg_success_10 ? _GEN_2215 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2361 = next_reg_vmEnable_10 ? _GEN_2345 : _GEN_2215; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_2410 = _T_846 ? _GEN_2361 : _GEN_2215; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire  _GEN_2468 = _T_393 ? _GEN_2410 : _GEN_2215; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire  _GEN_2598 = next_reg_success_10 ? _GEN_2468 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2614 = next_reg_vmEnable_10 ? _GEN_2598 : _GEN_2468; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_2663 = _T_848 ? _GEN_2614 : _GEN_2468; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire  _GEN_2721 = _T_413 ? _GEN_2663 : _GEN_2468; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2853 = next_reg_success_10 ? _GEN_2721 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2869 = next_reg_vmEnable_10 ? _GEN_2853 : _GEN_2721; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_2927 = _T_433 ? _GEN_2869 : _GEN_2721; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire  _GEN_3055 = next_reg_success_10 ? _GEN_2927 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_3071 = next_reg_vmEnable_10 ? _GEN_3055 : _GEN_2927; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_3120 = _T_846 ? _GEN_3071 : _GEN_2927; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire  _GEN_3178 = _T_452 ? _GEN_3120 : _GEN_2927; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire  _GEN_4871 = next_reg_success_10 ? _GEN_3178 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_4887 = next_reg_vmEnable_10 ? _GEN_4871 : _GEN_3178; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_4936 = _T_848 ? _GEN_4887 : _GEN_3178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire  _GEN_4994 = _T_818 ? _GEN_4936 : _GEN_3178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire  _GEN_5124 = next_reg_success_10 ? _GEN_4994 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5140 = next_reg_vmEnable_10 ? _GEN_5124 : _GEN_4994; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_5189 = _T_850 ? _GEN_5140 : _GEN_4994; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire  _GEN_5247 = _T_838 ? _GEN_5189 : _GEN_4994; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire  _GEN_5537 = next_reg_success_10 ? _GEN_5247 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5553 = next_reg_vmEnable_10 ? _GEN_5537 : _GEN_5247; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_5610 = _T_937 ? _GEN_5553 : _GEN_5247; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire  _GEN_5908 = next_reg_success_10 ? _GEN_5610 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5924 = next_reg_vmEnable_10 ? _GEN_5908 : _GEN_5610; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_5981 = _T_1005 ? _GEN_5924 : _GEN_5610; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire  _GEN_7827 = next_reg_success_10 ? _GEN_5981 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_7843 = next_reg_vmEnable_10 ? _GEN_7827 : _GEN_5981; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_7900 = _T_1308 ? _GEN_7843 : _GEN_5981; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire  _GEN_8198 = next_reg_success_10 ? _GEN_7900 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_8214 = next_reg_vmEnable_10 ? _GEN_8198 : _GEN_7900; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_8271 = _T_1376 ? _GEN_8214 : _GEN_7900; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire  exceptionVec_13 = io_valid & _GEN_8271; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_2 = exceptionVec_13 ? 6'hd : 6'h0; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _GEN_8404 = next_reg_permStore_10 & _GEN_8164; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 346:11 371:24]
  wire  success_8 = ~(next_reg_successLevel_10 == 2'h3) & _GEN_8404; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 335:37 376:22]
  wire  _GEN_3310 = success_8 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30 144:33]
  wire  _GEN_3326 = next_reg_vmEnable_10 & _GEN_3310; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_3353 = _T_472 & _GEN_3326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_3450 = success_8 ? _GEN_3353 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_3466 = next_reg_vmEnable_10 ? _GEN_3450 : _GEN_3353; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_3483 = _T_846 ? _GEN_3466 : _GEN_3353; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55]
  wire  _GEN_3511 = _T_547 ? _GEN_3483 : _GEN_3353; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire  _GEN_3610 = success_8 ? _GEN_3511 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_3626 = next_reg_vmEnable_10 ? _GEN_3610 : _GEN_3511; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_3643 = _T_848 ? _GEN_3626 : _GEN_3511; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55]
  wire  _GEN_3671 = _T_623 ? _GEN_3643 : _GEN_3511; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire  _GEN_5377 = success_8 ? _GEN_3671 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5393 = next_reg_vmEnable_10 ? _GEN_5377 : _GEN_3671; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_5410 = _T_850 ? _GEN_5393 : _GEN_3671; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55]
  wire  _GEN_5438 = _T_858 ? _GEN_5410 : _GEN_3671; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire  _GEN_5739 = success_8 ? _GEN_5438 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5755 = next_reg_vmEnable_10 ? _GEN_5739 : _GEN_5438; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_5778 = _T_944 ? _GEN_5755 : _GEN_5438; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24]
  wire  _GEN_6142 = success_8 ? _GEN_5778 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_6158 = next_reg_vmEnable_10 ? _GEN_6142 : _GEN_5778; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_6215 = _T_1014 ? _GEN_6158 : _GEN_5778; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22]
  wire  _GEN_8029 = success_8 ? _GEN_6215 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_8045 = next_reg_vmEnable_10 ? _GEN_8029 : _GEN_6215; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_8068 = _T_1315 ? _GEN_8045 : _GEN_6215; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24]
  wire  _GEN_8432 = success_8 ? _GEN_8068 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_8448 = next_reg_vmEnable_10 ? _GEN_8432 : _GEN_8068; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_8505 = _T_1385 ? _GEN_8448 : _GEN_8068; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22]
  wire  exceptionVec_15 = io_valid & _GEN_8505; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_3 = exceptionVec_15 ? 6'hf : _exceptionNO_T_2; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [4:0] _GEN_945 = _T_88 ? inst[24:20] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 20:24]
  wire [4:0] _GEN_1016 = _T_95 ? inst[24:20] : _GEN_945; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1087 = _T_102 ? inst[24:20] : _GEN_1016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1158 = _T_109 ? inst[24:20] : _GEN_1087; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1229 = _T_116 ? inst[24:20] : _GEN_1158; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1300 = _T_123 ? inst[24:20] : _GEN_1229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1371 = _T_762 ? inst[24:20] : _GEN_1300; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1442 = _T_769 ? inst[24:20] : _GEN_1371; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1513 = _T_144 ? inst[24:20] : _GEN_1442; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1584 = _T_776 ? inst[24:20] : _GEN_1513; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1861 = _T_207 ? inst[24:20] : _GEN_1584; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1886 = _T_234 ? inst[24:20] : _GEN_1861; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1911 = _T_261 ? inst[24:20] : _GEN_1886; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1936 = _T_290 ? inst[24:20] : _GEN_1911; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1961 = _T_317 ? inst[24:20] : _GEN_1936; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1986 = _T_346 ? inst[24:20] : _GEN_1961; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3330 = _T_472 ? inst[24:20] : _GEN_1986; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3490 = _T_547 ? inst[24:20] : _GEN_3330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3650 = _T_623 ? inst[24:20] : _GEN_3490; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4243 = _T_762 ? inst[24:20] : _GEN_3650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4314 = _T_769 ? inst[24:20] : _GEN_4243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4385 = _T_776 ? inst[24:20] : _GEN_4314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4456 = _T_783 ? inst[24:20] : _GEN_4385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4527 = _T_790 ? inst[24:20] : _GEN_4456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4598 = _T_797 ? inst[24:20] : _GEN_4527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4669 = _T_804 ? inst[24:20] : _GEN_4598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4740 = _T_811 ? inst[24:20] : _GEN_4669; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5417 = _T_858 ? inst[24:20] : _GEN_4740; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5760 = _T_944 ? inst[6:2] : _GEN_5417; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6237 = _T_1092 ? inst[6:2] : _GEN_5760; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_6245 = _T_1101 ? inst[6:2] : _GEN_6237; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7081 = _T_1248 ? inst[6:2] : _GEN_6245; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_7151 = _T_1260 ? inst[6:2] : _GEN_7081; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_8050 = _T_1315 ? inst[6:2] : _GEN_7151; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_8885 = _T_1475 ? inst[24:20] : _GEN_8050; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_8956 = _T_1482 ? inst[24:20] : _GEN_8885; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9027 = _T_1489 ? inst[24:20] : _GEN_8956; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9098 = _T_1496 ? inst[24:20] : _GEN_9027; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9169 = _T_1503 ? inst[24:20] : _GEN_9098; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9240 = _T_1510 ? inst[24:20] : _GEN_9169; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9311 = _T_1517 ? inst[24:20] : _GEN_9240; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9382 = _T_1524 ? inst[24:20] : _GEN_9311; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9453 = _T_1531 ? inst[24:20] : _GEN_9382; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9524 = _T_1538 ? inst[24:20] : _GEN_9453; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9595 = _T_1545 ? inst[24:20] : _GEN_9524; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9666 = _T_1552 ? inst[24:20] : _GEN_9595; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9737 = _T_1559 ? inst[24:20] : _GEN_9666; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] rs2 = io_valid ? _GEN_9737 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 20:24]
  wire  _GEN_2445 = _T_846 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2503 = _T_393 & _GEN_2445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire  _GEN_2698 = _T_848 ? _GEN_2503 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_2756 = _T_413 ? _GEN_2698 : _GEN_2503; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_3155 = _T_846 ? _GEN_2756 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_3213 = _T_452 ? _GEN_3155 : _GEN_2756; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire  _GEN_4971 = _T_848 ? _GEN_3213 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5029 = _T_818 ? _GEN_4971 : _GEN_3213; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire  _GEN_5224 = _T_850 ? _GEN_5029 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5282 = _T_838 ? _GEN_5224 : _GEN_5029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire  exceptionVec_4 = io_valid & _GEN_5282; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_4 = exceptionVec_4 ? 6'h4 : _exceptionNO_T_3; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _GEN_3515 = _T_547 & _GEN_2445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire  _GEN_3647 = _T_848 ? _GEN_3515 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_3675 = _T_623 ? _GEN_3647 : _GEN_3515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire  _GEN_5414 = _T_850 ? _GEN_3675 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_5442 = _T_858 ? _GEN_5414 : _GEN_3675; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire  exceptionVec_6 = io_valid & _GEN_5442; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_5 = exceptionVec_6 ? 6'h6 : _exceptionNO_T_4; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _T_710 = 2'h3 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42]
  wire  _GEN_3689 = 2'h1 == io_now_internal_privilegeMode ? 1'h0 : 2'h0 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_3693 = 2'h3 == io_now_internal_privilegeMode ? 1'h0 : _GEN_3689; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_3704 = _T_705 & _GEN_3693; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  exceptionVec_8 = io_valid & _GEN_3704; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_6 = exceptionVec_8 ? 6'h8 : _exceptionNO_T_5; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _GEN_3692 = 2'h3 == io_now_internal_privilegeMode ? 1'h0 : 2'h1 == io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_3703 = _T_705 & _GEN_3692; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  exceptionVec_9 = io_valid & _GEN_3703; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_7 = exceptionVec_9 ? 6'h9 : _exceptionNO_T_6; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  _GEN_3701 = _T_705 & _T_710; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  exceptionVec_11 = io_valid & _GEN_3701; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_8 = exceptionVec_11 ? 6'hb : _exceptionNO_T_7; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _GEN_880 = 5'h1 == rs2 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_881 = 5'h2 == rs2 ? io_now_reg_2 : _GEN_880; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_882 = 5'h3 == rs2 ? io_now_reg_3 : _GEN_881; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_883 = 5'h4 == rs2 ? io_now_reg_4 : _GEN_882; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_884 = 5'h5 == rs2 ? io_now_reg_5 : _GEN_883; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_885 = 5'h6 == rs2 ? io_now_reg_6 : _GEN_884; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_886 = 5'h7 == rs2 ? io_now_reg_7 : _GEN_885; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_887 = 5'h8 == rs2 ? io_now_reg_8 : _GEN_886; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_888 = 5'h9 == rs2 ? io_now_reg_9 : _GEN_887; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_889 = 5'ha == rs2 ? io_now_reg_10 : _GEN_888; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_890 = 5'hb == rs2 ? io_now_reg_11 : _GEN_889; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_891 = 5'hc == rs2 ? io_now_reg_12 : _GEN_890; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_892 = 5'hd == rs2 ? io_now_reg_13 : _GEN_891; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_893 = 5'he == rs2 ? io_now_reg_14 : _GEN_892; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_894 = 5'hf == rs2 ? io_now_reg_15 : _GEN_893; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_895 = 5'h10 == rs2 ? io_now_reg_16 : _GEN_894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_896 = 5'h11 == rs2 ? io_now_reg_17 : _GEN_895; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_897 = 5'h12 == rs2 ? io_now_reg_18 : _GEN_896; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_898 = 5'h13 == rs2 ? io_now_reg_19 : _GEN_897; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_899 = 5'h14 == rs2 ? io_now_reg_20 : _GEN_898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_900 = 5'h15 == rs2 ? io_now_reg_21 : _GEN_899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_901 = 5'h16 == rs2 ? io_now_reg_22 : _GEN_900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_902 = 5'h17 == rs2 ? io_now_reg_23 : _GEN_901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_903 = 5'h18 == rs2 ? io_now_reg_24 : _GEN_902; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_904 = 5'h19 == rs2 ? io_now_reg_25 : _GEN_903; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_905 = 5'h1a == rs2 ? io_now_reg_26 : _GEN_904; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_906 = 5'h1b == rs2 ? io_now_reg_27 : _GEN_905; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_907 = 5'h1c == rs2 ? io_now_reg_28 : _GEN_906; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_908 = 5'h1d == rs2 ? io_now_reg_29 : _GEN_907; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_909 = 5'h1e == rs2 ? io_now_reg_30 : _GEN_908; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [63:0] _GEN_910 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_909; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{62,62}]
  wire [1:0] _T_357 = io_now_csr_misa[2] ? 2'h1 : 2'h2; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 134:62]
  wire [63:0] _T_359 = io_now_pc + imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:49]
  wire  _T_365 = _T_359[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_363 = _T_359[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_361 = ~_T_359[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_367 = 2'h1 == _T_357 ? _T_361 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_369 = 2'h2 == _T_357 ? _T_363 : _T_367; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_371 = 2'h3 == _T_357 ? _T_365 : _T_369; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire [63:0] _T_325 = 5'h1f == rs1 ? io_now_reg_31 : _GEN_100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:25]
  wire [63:0] _T_326 = 5'h1f == rs2 ? io_now_reg_31 : _GEN_909; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:48]
  wire  _T_298 = _GEN_101 < _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:25]
  wire  _T_271 = $signed(_T_325) < $signed(_T_326); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:32]
  wire [63:0] _T_193 = {_T_844[63:1],1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:43]
  wire  _T_199 = _T_193[2:0] == 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 128:32]
  wire  _T_197 = _T_193[1:0] == 2'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 127:32]
  wire  _T_195 = ~_T_193[0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 126:29]
  wire  _T_201 = 2'h1 == _T_357 ? _T_195 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_203 = 2'h2 == _T_357 ? _T_197 : _T_201; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _T_205 = 2'h3 == _T_357 ? _T_199 : _T_203; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 123:29]
  wire  _GEN_1688 = _T_371 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30 144:33]
  wire  _GEN_1733 = _T_158 & _GEN_1688; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_1802 = _T_205 ? _GEN_1733 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1846 = _T_182 ? _GEN_1802 : _GEN_1733; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire  _GEN_1851 = _T_371 ? _GEN_1846 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1856 = _GEN_101 == _GEN_910 ? _GEN_1851 : _GEN_1846; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire  _GEN_1871 = _T_207 ? _GEN_1856 : _GEN_1846; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire  _GEN_1876 = _T_371 ? _GEN_1871 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1881 = _GEN_101 != _GEN_910 ? _GEN_1876 : _GEN_1871; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire  _GEN_1896 = _T_234 ? _GEN_1881 : _GEN_1871; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire  _GEN_1901 = _T_371 ? _GEN_1896 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1906 = $signed(_T_325) < $signed(_T_326) ? _GEN_1901 : _GEN_1896; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire  _GEN_1921 = _T_261 ? _GEN_1906 : _GEN_1896; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire  _GEN_1926 = _T_371 ? _GEN_1921 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1931 = _GEN_101 < _GEN_910 ? _GEN_1926 : _GEN_1921; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire  _GEN_1946 = _T_290 ? _GEN_1931 : _GEN_1921; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire  _GEN_1951 = _T_371 ? _GEN_1946 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1956 = $signed(_T_325) >= $signed(_T_326) ? _GEN_1951 : _GEN_1946; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire  _GEN_1971 = _T_317 ? _GEN_1956 : _GEN_1946; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire  _GEN_1976 = _T_371 ? _GEN_1971 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_1981 = _GEN_101 >= _GEN_910 ? _GEN_1976 : _GEN_1971; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire  _GEN_1996 = _T_346 ? _GEN_1981 : _GEN_1971; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire  exceptionVec_0 = io_valid & _GEN_1996; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_9 = exceptionVec_0 ? 6'h0 : _exceptionNO_T_8; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _T_1466 = inst & 32'hfc63; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1467 = 32'h9c01 == _T_1466; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1459 = 32'h9c21 == _T_1466; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1290 = 32'h8c01 == _T_1466; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1282 = 32'h8c21 == _T_1466; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1274 = 32'h8c41 == _T_1466; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1266 = 32'h8c61 == _T_1466; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_1182 = inst[12:5] != 8'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 23:96]
  wire  _T_1183 = 32'h0 == _T_1375 & _T_1182; // @[src/main/scala/rvspeccore/core/spec/RVInsts.scala 11:45]
  wire  _GEN_134 = _T_26 ? 1'h0 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 125:24 128:24]
  wire  _GEN_205 = _T_32 ? 1'h0 : _GEN_134; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_276 = _T_38 ? 1'h0 : _GEN_205; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_347 = _T_44 ? 1'h0 : _GEN_276; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_418 = _T_50 ? 1'h0 : _GEN_347; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_489 = _T_56 ? 1'h0 : _GEN_418; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_560 = _T_726 ? 1'h0 : _GEN_489; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_631 = _T_732 ? 1'h0 : _GEN_560; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_702 = _T_738 ? 1'h0 : _GEN_631; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_773 = _T_80 ? 1'h0 : _GEN_702; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_842 = _T_84 ? 1'h0 : _GEN_773; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_943 = _T_88 ? 1'h0 : _GEN_842; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1014 = _T_95 ? 1'h0 : _GEN_943; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1085 = _T_102 ? 1'h0 : _GEN_1014; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1156 = _T_109 ? 1'h0 : _GEN_1085; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1227 = _T_116 ? 1'h0 : _GEN_1156; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1298 = _T_123 ? 1'h0 : _GEN_1227; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1369 = _T_762 ? 1'h0 : _GEN_1298; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1440 = _T_769 ? 1'h0 : _GEN_1369; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1511 = _T_144 ? 1'h0 : _GEN_1440; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1582 = _T_776 ? 1'h0 : _GEN_1511; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1690 = _T_158 ? 1'h0 : _GEN_1582; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1804 = _T_182 ? 1'h0 : _GEN_1690; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1858 = _T_207 ? 1'h0 : _GEN_1804; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1883 = _T_234 ? 1'h0 : _GEN_1858; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1908 = _T_261 ? 1'h0 : _GEN_1883; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1933 = _T_290 ? 1'h0 : _GEN_1908; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1958 = _T_317 ? 1'h0 : _GEN_1933; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_1983 = _T_346 ? 1'h0 : _GEN_1958; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2193 = _T_373 ? 1'h0 : _GEN_1983; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2446 = _T_393 ? 1'h0 : _GEN_2193; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2699 = _T_413 ? 1'h0 : _GEN_2446; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_2903 = _T_433 ? 1'h0 : _GEN_2699; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3156 = _T_452 ? 1'h0 : _GEN_2903; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3328 = _T_472 ? 1'h0 : _GEN_3156; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3488 = _T_547 ? 1'h0 : _GEN_3328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3648 = _T_623 ? 1'h0 : _GEN_3488; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3676 = _T_699 ? 1'h0 : _GEN_3648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3694 = _T_705 ? 1'h0 : _GEN_3676; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3705 = _T_714 ? 1'h0 : _GEN_3694; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3744 = _T_720 ? 1'h0 : _GEN_3705; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3815 = _T_726 ? 1'h0 : _GEN_3744; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3886 = _T_732 ? 1'h0 : _GEN_3815; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_3957 = _T_738 ? 1'h0 : _GEN_3886; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4028 = _T_744 ? 1'h0 : _GEN_3957; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4099 = _T_750 ? 1'h0 : _GEN_4028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4170 = _T_756 ? 1'h0 : _GEN_4099; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4241 = _T_762 ? 1'h0 : _GEN_4170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4312 = _T_769 ? 1'h0 : _GEN_4241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4383 = _T_776 ? 1'h0 : _GEN_4312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4454 = _T_783 ? 1'h0 : _GEN_4383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4525 = _T_790 ? 1'h0 : _GEN_4454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4596 = _T_797 ? 1'h0 : _GEN_4525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4667 = _T_804 ? 1'h0 : _GEN_4596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4738 = _T_811 ? 1'h0 : _GEN_4667; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_4972 = _T_818 ? 1'h0 : _GEN_4738; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5225 = _T_838 ? 1'h0 : _GEN_4972; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5415 = _T_858 ? 1'h0 : _GEN_5225; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5587 = _T_937 ? 1'h0 : _GEN_5415; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5757 = _T_944 ? 1'h0 : _GEN_5587; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_5958 = _T_1005 ? 1'h0 : _GEN_5757; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6192 = _T_1014 ? 1'h0 : _GEN_5958; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6219 = _T_1078 ? 1'h0 : _GEN_6192; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 160:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6234 = _T_1092 ? 1'h0 : _GEN_6219; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6242 = _T_1101 ? 1'h0 : _GEN_6234; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6285 = _T_1107 ? 1'h0 : _GEN_6242; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6329 = _T_1116 ? 1'h0 : _GEN_6285; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6371 = _T_1128 ? 1'h0 : _GEN_6329; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6443 = _T_1146 ? 1'h0 : _GEN_6371; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6546 = _T_1161 ? 1'h0 : _GEN_6443; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6585 = _T_1173 ? 1'h0 : _GEN_6546; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 220:28 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6625 = _T_1183 ? 1'h0 : _GEN_6585; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6694 = _T_1199 ? 1'h0 : _GEN_6625; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6798 = _T_1212 ? 1'h0 : _GEN_6694; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_6902 = _T_1226 ? 1'h0 : _GEN_6798; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_7006 = _T_1234 ? 1'h0 : _GEN_6902; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_7078 = _T_1248 ? 1'h0 : _GEN_7006; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_7148 = _T_1260 ? 1'h0 : _GEN_7078; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_7282 = _T_1266 ? 1'h0 : _GEN_7148; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_7417 = _T_1274 ? 1'h0 : _GEN_7282; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_7552 = _T_1282 ? 1'h0 : _GEN_7417; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_7687 = _T_1290 ? 1'h0 : _GEN_7552; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_7726 = _T_1298 ? 1'h0 : _GEN_7687; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 259:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_7877 = _T_1308 ? 1'h0 : _GEN_7726; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_8047 = _T_1315 ? 1'h0 : _GEN_7877; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_8248 = _T_1376 ? 1'h0 : _GEN_8047; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_8482 = _T_1385 ? 1'h0 : _GEN_8248; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_8541 = _T_1452 ? 1'h0 : _GEN_8482; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_8677 = _T_1459 ? 1'h0 : _GEN_8541; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_8812 = _T_1467 ? 1'h0 : _GEN_8677; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_8883 = _T_1475 ? 1'h0 : _GEN_8812; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_8954 = _T_1482 ? 1'h0 : _GEN_8883; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_9025 = _T_1489 ? 1'h0 : _GEN_8954; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_9096 = _T_1496 ? 1'h0 : _GEN_9025; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_9167 = _T_1503 ? 1'h0 : _GEN_9096; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_9238 = _T_1510 ? 1'h0 : _GEN_9167; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_9309 = _T_1517 ? 1'h0 : _GEN_9238; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_9380 = _T_1524 ? 1'h0 : _GEN_9309; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_9451 = _T_1531 ? 1'h0 : _GEN_9380; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_9522 = _T_1538 ? 1'h0 : _GEN_9451; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_9593 = _T_1545 ? 1'h0 : _GEN_9522; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_9664 = _T_1552 ? 1'h0 : _GEN_9593; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_9735 = _T_1559 ? 1'h0 : _GEN_9664; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_9785 = _T_1566 ? 1'h0 : _GEN_9735; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_9806 = _T_1573 ? 1'h0 : _GEN_9785; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_9820 = _T_1580 ? 1'h0 : _GEN_9806; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_9827 = _T_1586 ? 1'h0 : _GEN_9820; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_9974 = _T_1592 ? 1'h0 : _GEN_9827; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_10154 = _T_1625 ? 1'h0 : _GEN_9974; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_10334 = _T_1667 ? 1'h0 : _GEN_10154; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_10526 = _T_1709 ? 1'h0 : _GEN_10334; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_10706 = _T_1743 ? 1'h0 : _GEN_10526; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  _GEN_10886 = _T_1786 ? 1'h0 : _GEN_10706; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 128:24]
  wire  illegalInstruction = io_valid & _GEN_10886; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 119:36]
  wire [11:0] _GEN_9981 = _T_1592 ? imm[11:0] : 12'h0; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 56:13 82:23 53:25]
  wire [11:0] _GEN_10161 = _T_1625 ? imm[11:0] : _GEN_9981; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 56:13 93:23]
  wire [11:0] _GEN_10341 = _T_1667 ? imm[11:0] : _GEN_10161; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23 56:13]
  wire [11:0] _GEN_10533 = _T_1709 ? imm[11:0] : _GEN_10341; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24 56:13]
  wire [11:0] _GEN_10713 = _T_1743 ? imm[11:0] : _GEN_10533; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24 56:13]
  wire [11:0] _GEN_10893 = _T_1786 ? imm[11:0] : _GEN_10713; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24 56:13]
  wire [11:0] csrAddr = io_valid ? _GEN_10893 : 12'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 53:25]
  wire  isIllegalWrite_5 = csrAddr[11:10] == 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:39]
  wire  _T_1793 = ~isIllegalWrite_5; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:12]
  wire  _T_1794 = rs1 != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:18]
  wire  _has_T_431 = 12'h343 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_429 = 12'h342 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_427 = 12'h341 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_425 = 12'h304 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_423 = 12'h344 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_421 = 12'h306 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_419 = 12'h305 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_417 = 12'h340 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_415 = 12'h300 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_413 = 12'hf14 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_411 = 12'hf13 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_409 = 12'hf12 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_407 = 12'hf11 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  _has_T_405 = 12'h301 == csrAddr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  has_15 = 12'h343 == csrAddr | (12'h342 == csrAddr | (12'h341 == csrAddr | (12'h304 == csrAddr | (12'h344 ==
    csrAddr | (12'h306 == csrAddr | (12'h305 == csrAddr | (12'h340 == csrAddr | (12'h300 == csrAddr | (12'hf14 ==
    csrAddr | (12'hf13 == csrAddr | (12'hf12 == csrAddr | (12'hf11 == csrAddr | 12'h301 == csrAddr)))))))))))); // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 61:45]
  wire  isIllegalMode_5 = io_now_internal_privilegeMode < csrAddr[9:8]; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 72:53]
  wire  isIllegalAccess_5 = isIllegalMode_5 | isIllegalWrite_5; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 74:41]
  wire  _T_1748 = _GEN_101 == 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:39]
  wire  isIllegalWrite_4 = isIllegalWrite_5 & ~_T_1748; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 71:51]
  wire  _T_1751 = ~isIllegalWrite_4; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:12]
  wire  isIllegalAccess_4 = isIllegalMode_5 | isIllegalWrite_4; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 74:41]
  wire  illegalSret = io_now_internal_privilegeMode < 2'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 118:55]
  wire  mstatusOld_tsr = io_now_csr_mstatus[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 111:55]
  wire  illegalSModeSret = io_now_internal_privilegeMode == 2'h1 & mstatusOld_tsr; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 119:65]
  wire  _T_1571 = illegalSret | illegalSModeSret; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:22]
  wire  _GEN_9792 = _T_1566 & _T_1571; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire  _GEN_9804 = io_now_internal_privilegeMode == 2'h3 ? _GEN_9792 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 88:48 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_9818 = _T_1573 ? _GEN_9804 : _GEN_9792; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire  _GEN_9834 = isIllegalAccess_5 | ~has_15 | _GEN_9818; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_9928 = has_15 ? _GEN_9834 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_9972 = _T_1793 ? _GEN_9928 : _GEN_9834; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire  _GEN_9982 = _T_1592 ? _GEN_9972 : _GEN_9818; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire  _GEN_10026 = isIllegalAccess_4 | ~has_15 | _GEN_9982; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_10096 = has_15 ? _GEN_10026 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_10108 = _T_1794 ? _GEN_10096 : _GEN_10026; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire  _GEN_10152 = _T_1751 ? _GEN_10108 : _GEN_10026; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire  _GEN_10162 = _T_1625 ? _GEN_10152 : _GEN_9982; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire  _GEN_10206 = isIllegalAccess_5 | ~has_15 | _GEN_10162; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_10276 = has_15 ? _GEN_10206 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_10288 = _T_1794 ? _GEN_10276 : _GEN_10206; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire  _GEN_10332 = _T_1793 ? _GEN_10288 : _GEN_10206; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire  _GEN_10342 = _T_1667 ? _GEN_10332 : _GEN_10162; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire  _GEN_10386 = isIllegalAccess_5 | ~has_15 | _GEN_10342; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_10480 = has_15 ? _GEN_10386 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_10524 = _T_1793 ? _GEN_10480 : _GEN_10386; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire  _GEN_10534 = _T_1709 ? _GEN_10524 : _GEN_10342; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire  _GEN_10578 = isIllegalAccess_4 | ~has_15 | _GEN_10534; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_10648 = has_15 ? _GEN_10578 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_10660 = _T_1794 ? _GEN_10648 : _GEN_10578; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire  _GEN_10704 = ~isIllegalWrite_4 ? _GEN_10660 : _GEN_10578; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire  _GEN_10714 = _T_1743 ? _GEN_10704 : _GEN_10534; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire  _GEN_10758 = isIllegalAccess_5 | ~has_15 | _GEN_10714; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_10828 = has_15 ? _GEN_10758 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 144:33]
  wire  _GEN_10840 = rs1 != 5'h0 ? _GEN_10828 : _GEN_10758; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire  _GEN_10884 = ~isIllegalWrite_5 ? _GEN_10840 : _GEN_10758; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire  _GEN_10894 = _T_1786 ? _GEN_10884 : _GEN_10714; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire  _GEN_10939 = illegalInstruction | _GEN_10894; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 133:30 144:33]
  wire  exceptionVec_2 = io_valid & _GEN_10939; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_10 = exceptionVec_2 ? 6'h2 : _exceptionNO_T_9; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  exceptionVec_12 = io_valid & vmEnable; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] _exceptionNO_T_12 = exceptionVec_12 ? 6'hc : _exceptionNO_T_10; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  exceptionVec_3 = io_valid & _T_699; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 122:30]
  wire [5:0] exceptionNO = exceptionVec_3 ? 6'h3 : _exceptionNO_T_12; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [4:0] _GEN_138 = _T_26 ? inst[11:7] : 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 17:24]
  wire [4:0] _GEN_209 = _T_32 ? inst[11:7] : _GEN_138; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_280 = _T_38 ? inst[11:7] : _GEN_209; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_351 = _T_44 ? inst[11:7] : _GEN_280; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_422 = _T_50 ? inst[11:7] : _GEN_351; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_493 = _T_56 ? inst[11:7] : _GEN_422; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_564 = _T_726 ? inst[11:7] : _GEN_493; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_635 = _T_732 ? inst[11:7] : _GEN_564; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_706 = _T_738 ? inst[11:7] : _GEN_635; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_775 = _T_80 ? inst[11:7] : _GEN_706; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_844 = _T_84 ? inst[11:7] : _GEN_775; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_948 = _T_88 ? inst[11:7] : _GEN_844; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1019 = _T_95 ? inst[11:7] : _GEN_948; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1090 = _T_102 ? inst[11:7] : _GEN_1019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1161 = _T_109 ? inst[11:7] : _GEN_1090; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1232 = _T_116 ? inst[11:7] : _GEN_1161; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1303 = _T_123 ? inst[11:7] : _GEN_1232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1374 = _T_762 ? inst[11:7] : _GEN_1303; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1445 = _T_769 ? inst[11:7] : _GEN_1374; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1516 = _T_144 ? inst[11:7] : _GEN_1445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1587 = _T_776 ? inst[11:7] : _GEN_1516; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1695 = _T_158 ? inst[11:7] : _GEN_1587; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_1808 = _T_182 ? inst[11:7] : _GEN_1695; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2197 = _T_373 ? inst[11:7] : _GEN_1808; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2450 = _T_393 ? inst[11:7] : _GEN_2197; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2703 = _T_413 ? inst[11:7] : _GEN_2450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_2907 = _T_433 ? inst[11:7] : _GEN_2703; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3160 = _T_452 ? inst[11:7] : _GEN_2907; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3680 = _T_699 ? inst[11:7] : _GEN_3160; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3698 = _T_705 ? inst[11:7] : _GEN_3680; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3709 = _T_714 ? inst[11:7] : _GEN_3698; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 360:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3748 = _T_720 ? inst[11:7] : _GEN_3709; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3819 = _T_726 ? inst[11:7] : _GEN_3748; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3890 = _T_732 ? inst[11:7] : _GEN_3819; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_3961 = _T_738 ? inst[11:7] : _GEN_3890; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4032 = _T_744 ? inst[11:7] : _GEN_3961; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4103 = _T_750 ? inst[11:7] : _GEN_4032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4174 = _T_756 ? inst[11:7] : _GEN_4103; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4246 = _T_762 ? inst[11:7] : _GEN_4174; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4317 = _T_769 ? inst[11:7] : _GEN_4246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4388 = _T_776 ? inst[11:7] : _GEN_4317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4459 = _T_783 ? inst[11:7] : _GEN_4388; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4530 = _T_790 ? inst[11:7] : _GEN_4459; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4601 = _T_797 ? inst[11:7] : _GEN_4530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4672 = _T_804 ? inst[11:7] : _GEN_4601; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4743 = _T_811 ? inst[11:7] : _GEN_4672; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_4976 = _T_818 ? inst[11:7] : _GEN_4743; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5229 = _T_838 ? inst[11:7] : _GEN_4976; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_5593 = _T_937 ? rs1 : _GEN_5229; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 138:24]
  wire [4:0] _GEN_6239 = _T_1092 ? rs1 : _GEN_5593; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 112:110 173:22]
  wire [4:0] _GEN_6247 = _T_1101 ? rs1 : _GEN_6239; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 112:110 179:24]
  wire [4:0] _GEN_6377 = _T_1128 ? rs1 : _GEN_6247; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 204:22]
  wire [4:0] _GEN_6449 = _T_1146 ? rs1 : _GEN_6377; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 209:23]
  wire [4:0] _GEN_6552 = _T_1161 ? rs1 : _GEN_6449; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 215:24]
  wire [4:0] _GEN_6591 = _T_1173 ? rs1 : _GEN_6552; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 220:28]
  wire [4:0] _GEN_6700 = _T_1199 ? rs1 : _GEN_6591; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 230:24]
  wire [4:0] _GEN_7083 = _T_1248 ? rs1 : _GEN_6700; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 112:110 251:23]
  wire [4:0] _GEN_7153 = _T_1260 ? rs1 : _GEN_7083; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 112:110 252:23]
  wire [4:0] _GEN_7732 = _T_1298 ? rs1 : _GEN_7153; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 259:23]
  wire [4:0] _GEN_7883 = _T_1308 ? rs1 : _GEN_7732; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 267:24]
  wire [4:0] _GEN_8547 = _T_1452 ? rs1 : _GEN_7883; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 113:110 290:25]
  wire [4:0] _GEN_8888 = _T_1475 ? inst[11:7] : _GEN_8547; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_8959 = _T_1482 ? inst[11:7] : _GEN_8888; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9030 = _T_1489 ? inst[11:7] : _GEN_8959; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9101 = _T_1496 ? inst[11:7] : _GEN_9030; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9172 = _T_1503 ? inst[11:7] : _GEN_9101; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9243 = _T_1510 ? inst[11:7] : _GEN_9172; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9314 = _T_1517 ? inst[11:7] : _GEN_9243; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9385 = _T_1524 ? inst[11:7] : _GEN_9314; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9456 = _T_1531 ? inst[11:7] : _GEN_9385; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9527 = _T_1538 ? inst[11:7] : _GEN_9456; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9598 = _T_1545 ? inst[11:7] : _GEN_9527; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9669 = _T_1552 ? inst[11:7] : _GEN_9598; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9740 = _T_1559 ? inst[11:7] : _GEN_9669; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9789 = _T_1566 ? inst[11:7] : _GEN_9740; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9810 = _T_1573 ? inst[11:7] : _GEN_9789; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9824 = _T_1580 ? inst[11:7] : _GEN_9810; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 62:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9831 = _T_1586 ? inst[11:7] : _GEN_9824; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 63:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_9978 = _T_1592 ? inst[11:7] : _GEN_9831; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_10158 = _T_1625 ? inst[11:7] : _GEN_9978; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_10338 = _T_1667 ? inst[11:7] : _GEN_10158; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_10530 = _T_1709 ? inst[11:7] : _GEN_10338; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_10710 = _T_1743 ? inst[11:7] : _GEN_10530; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] _GEN_10890 = _T_1786 ? inst[11:7] : _GEN_10710; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [4:0] rd = io_valid ? _GEN_10890 : 5'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CommonDecode.scala 17:24]
  wire [63:0] _GEN_103 = 5'h1 == rd ? _T_844 : io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_104 = 5'h2 == rd ? _T_844 : io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_105 = 5'h3 == rd ? _T_844 : io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_106 = 5'h4 == rd ? _T_844 : io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_107 = 5'h5 == rd ? _T_844 : io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_108 = 5'h6 == rd ? _T_844 : io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_109 = 5'h7 == rd ? _T_844 : io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_110 = 5'h8 == rd ? _T_844 : io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_111 = 5'h9 == rd ? _T_844 : io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_112 = 5'ha == rd ? _T_844 : io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_113 = 5'hb == rd ? _T_844 : io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_114 = 5'hc == rd ? _T_844 : io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_115 = 5'hd == rd ? _T_844 : io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_116 = 5'he == rd ? _T_844 : io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_117 = 5'hf == rd ? _T_844 : io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_118 = 5'h10 == rd ? _T_844 : io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_119 = 5'h11 == rd ? _T_844 : io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_120 = 5'h12 == rd ? _T_844 : io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_121 = 5'h13 == rd ? _T_844 : io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_122 = 5'h14 == rd ? _T_844 : io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_123 = 5'h15 == rd ? _T_844 : io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_124 = 5'h16 == rd ? _T_844 : io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_125 = 5'h17 == rd ? _T_844 : io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_126 = 5'h18 == rd ? _T_844 : io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_127 = 5'h19 == rd ? _T_844 : io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_128 = 5'h1a == rd ? _T_844 : io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_129 = 5'h1b == rd ? _T_844 : io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_130 = 5'h1c == rd ? _T_844 : io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_131 = 5'h1d == rd ? _T_844 : io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_132 = 5'h1e == rd ? _T_844 : io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_133 = 5'h1f == rd ? _T_844 : io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:{47,47}]
  wire [63:0] _GEN_142 = _T_26 ? _GEN_103 : io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_143 = _T_26 ? _GEN_104 : io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_144 = _T_26 ? _GEN_105 : io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_145 = _T_26 ? _GEN_106 : io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_146 = _T_26 ? _GEN_107 : io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_147 = _T_26 ? _GEN_108 : io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_148 = _T_26 ? _GEN_109 : io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_149 = _T_26 ? _GEN_110 : io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_150 = _T_26 ? _GEN_111 : io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_151 = _T_26 ? _GEN_112 : io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_152 = _T_26 ? _GEN_113 : io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_153 = _T_26 ? _GEN_114 : io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_154 = _T_26 ? _GEN_115 : io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_155 = _T_26 ? _GEN_116 : io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_156 = _T_26 ? _GEN_117 : io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_157 = _T_26 ? _GEN_118 : io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_158 = _T_26 ? _GEN_119 : io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_159 = _T_26 ? _GEN_120 : io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_160 = _T_26 ? _GEN_121 : io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_161 = _T_26 ? _GEN_122 : io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_162 = _T_26 ? _GEN_123 : io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_163 = _T_26 ? _GEN_124 : io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_164 = _T_26 ? _GEN_125 : io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_165 = _T_26 ? _GEN_126 : io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_166 = _T_26 ? _GEN_127 : io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_167 = _T_26 ? _GEN_128 : io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_168 = _T_26 ? _GEN_129 : io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_169 = _T_26 ? _GEN_130 : io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_170 = _T_26 ? _GEN_131 : io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_171 = _T_26 ? _GEN_132 : io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _GEN_172 = _T_26 ? _GEN_133 : io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 151:23]
  wire [63:0] _next_reg_T_3 = io_valid ? _GEN_10892 : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:80]
  wire [63:0] _next_reg_rd_0 = {{63'd0}, $signed(_T_325) < $signed(_next_reg_T_3)}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_174 = 5'h1 == rd ? _next_reg_rd_0 : _GEN_142; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_175 = 5'h2 == rd ? _next_reg_rd_0 : _GEN_143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_176 = 5'h3 == rd ? _next_reg_rd_0 : _GEN_144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_177 = 5'h4 == rd ? _next_reg_rd_0 : _GEN_145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_178 = 5'h5 == rd ? _next_reg_rd_0 : _GEN_146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_179 = 5'h6 == rd ? _next_reg_rd_0 : _GEN_147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_180 = 5'h7 == rd ? _next_reg_rd_0 : _GEN_148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_181 = 5'h8 == rd ? _next_reg_rd_0 : _GEN_149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_182 = 5'h9 == rd ? _next_reg_rd_0 : _GEN_150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_183 = 5'ha == rd ? _next_reg_rd_0 : _GEN_151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_184 = 5'hb == rd ? _next_reg_rd_0 : _GEN_152; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_185 = 5'hc == rd ? _next_reg_rd_0 : _GEN_153; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_186 = 5'hd == rd ? _next_reg_rd_0 : _GEN_154; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_187 = 5'he == rd ? _next_reg_rd_0 : _GEN_155; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_188 = 5'hf == rd ? _next_reg_rd_0 : _GEN_156; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_189 = 5'h10 == rd ? _next_reg_rd_0 : _GEN_157; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_190 = 5'h11 == rd ? _next_reg_rd_0 : _GEN_158; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_191 = 5'h12 == rd ? _next_reg_rd_0 : _GEN_159; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_192 = 5'h13 == rd ? _next_reg_rd_0 : _GEN_160; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_193 = 5'h14 == rd ? _next_reg_rd_0 : _GEN_161; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_194 = 5'h15 == rd ? _next_reg_rd_0 : _GEN_162; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_195 = 5'h16 == rd ? _next_reg_rd_0 : _GEN_163; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_196 = 5'h17 == rd ? _next_reg_rd_0 : _GEN_164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_197 = 5'h18 == rd ? _next_reg_rd_0 : _GEN_165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_198 = 5'h19 == rd ? _next_reg_rd_0 : _GEN_166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_199 = 5'h1a == rd ? _next_reg_rd_0 : _GEN_167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_200 = 5'h1b == rd ? _next_reg_rd_0 : _GEN_168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_201 = 5'h1c == rd ? _next_reg_rd_0 : _GEN_169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_202 = 5'h1d == rd ? _next_reg_rd_0 : _GEN_170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_203 = 5'h1e == rd ? _next_reg_rd_0 : _GEN_171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_204 = 5'h1f == rd ? _next_reg_rd_0 : _GEN_172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:{47,47}]
  wire [63:0] _GEN_213 = _T_32 ? _GEN_174 : _GEN_142; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_214 = _T_32 ? _GEN_175 : _GEN_143; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_215 = _T_32 ? _GEN_176 : _GEN_144; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_216 = _T_32 ? _GEN_177 : _GEN_145; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_217 = _T_32 ? _GEN_178 : _GEN_146; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_218 = _T_32 ? _GEN_179 : _GEN_147; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_219 = _T_32 ? _GEN_180 : _GEN_148; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_220 = _T_32 ? _GEN_181 : _GEN_149; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_221 = _T_32 ? _GEN_182 : _GEN_150; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_222 = _T_32 ? _GEN_183 : _GEN_151; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_223 = _T_32 ? _GEN_184 : _GEN_152; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_224 = _T_32 ? _GEN_185 : _GEN_153; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_225 = _T_32 ? _GEN_186 : _GEN_154; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_226 = _T_32 ? _GEN_187 : _GEN_155; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_227 = _T_32 ? _GEN_188 : _GEN_156; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_228 = _T_32 ? _GEN_189 : _GEN_157; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_229 = _T_32 ? _GEN_190 : _GEN_158; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_230 = _T_32 ? _GEN_191 : _GEN_159; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_231 = _T_32 ? _GEN_192 : _GEN_160; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_232 = _T_32 ? _GEN_193 : _GEN_161; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_233 = _T_32 ? _GEN_194 : _GEN_162; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_234 = _T_32 ? _GEN_195 : _GEN_163; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_235 = _T_32 ? _GEN_196 : _GEN_164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_236 = _T_32 ? _GEN_197 : _GEN_165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_237 = _T_32 ? _GEN_198 : _GEN_166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_238 = _T_32 ? _GEN_199 : _GEN_167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_239 = _T_32 ? _GEN_200 : _GEN_168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_240 = _T_32 ? _GEN_201 : _GEN_169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_241 = _T_32 ? _GEN_202 : _GEN_170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_242 = _T_32 ? _GEN_203 : _GEN_171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _GEN_243 = _T_32 ? _GEN_204 : _GEN_172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 152:23]
  wire [63:0] _next_reg_rd_1 = {{63'd0}, _GEN_101 < imm}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_245 = 5'h1 == rd ? _next_reg_rd_1 : _GEN_213; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_246 = 5'h2 == rd ? _next_reg_rd_1 : _GEN_214; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_247 = 5'h3 == rd ? _next_reg_rd_1 : _GEN_215; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_248 = 5'h4 == rd ? _next_reg_rd_1 : _GEN_216; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_249 = 5'h5 == rd ? _next_reg_rd_1 : _GEN_217; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_250 = 5'h6 == rd ? _next_reg_rd_1 : _GEN_218; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_251 = 5'h7 == rd ? _next_reg_rd_1 : _GEN_219; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_252 = 5'h8 == rd ? _next_reg_rd_1 : _GEN_220; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_253 = 5'h9 == rd ? _next_reg_rd_1 : _GEN_221; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_254 = 5'ha == rd ? _next_reg_rd_1 : _GEN_222; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_255 = 5'hb == rd ? _next_reg_rd_1 : _GEN_223; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_256 = 5'hc == rd ? _next_reg_rd_1 : _GEN_224; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_257 = 5'hd == rd ? _next_reg_rd_1 : _GEN_225; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_258 = 5'he == rd ? _next_reg_rd_1 : _GEN_226; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_259 = 5'hf == rd ? _next_reg_rd_1 : _GEN_227; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_260 = 5'h10 == rd ? _next_reg_rd_1 : _GEN_228; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_261 = 5'h11 == rd ? _next_reg_rd_1 : _GEN_229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_262 = 5'h12 == rd ? _next_reg_rd_1 : _GEN_230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_263 = 5'h13 == rd ? _next_reg_rd_1 : _GEN_231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_264 = 5'h14 == rd ? _next_reg_rd_1 : _GEN_232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_265 = 5'h15 == rd ? _next_reg_rd_1 : _GEN_233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_266 = 5'h16 == rd ? _next_reg_rd_1 : _GEN_234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_267 = 5'h17 == rd ? _next_reg_rd_1 : _GEN_235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_268 = 5'h18 == rd ? _next_reg_rd_1 : _GEN_236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_269 = 5'h19 == rd ? _next_reg_rd_1 : _GEN_237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_270 = 5'h1a == rd ? _next_reg_rd_1 : _GEN_238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_271 = 5'h1b == rd ? _next_reg_rd_1 : _GEN_239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_272 = 5'h1c == rd ? _next_reg_rd_1 : _GEN_240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_273 = 5'h1d == rd ? _next_reg_rd_1 : _GEN_241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_274 = 5'h1e == rd ? _next_reg_rd_1 : _GEN_242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_275 = 5'h1f == rd ? _next_reg_rd_1 : _GEN_243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:{47,47}]
  wire [63:0] _GEN_284 = _T_38 ? _GEN_245 : _GEN_213; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_285 = _T_38 ? _GEN_246 : _GEN_214; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_286 = _T_38 ? _GEN_247 : _GEN_215; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_287 = _T_38 ? _GEN_248 : _GEN_216; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_288 = _T_38 ? _GEN_249 : _GEN_217; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_289 = _T_38 ? _GEN_250 : _GEN_218; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_290 = _T_38 ? _GEN_251 : _GEN_219; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_291 = _T_38 ? _GEN_252 : _GEN_220; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_292 = _T_38 ? _GEN_253 : _GEN_221; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_293 = _T_38 ? _GEN_254 : _GEN_222; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_294 = _T_38 ? _GEN_255 : _GEN_223; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_295 = _T_38 ? _GEN_256 : _GEN_224; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_296 = _T_38 ? _GEN_257 : _GEN_225; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_297 = _T_38 ? _GEN_258 : _GEN_226; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_298 = _T_38 ? _GEN_259 : _GEN_227; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_299 = _T_38 ? _GEN_260 : _GEN_228; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_300 = _T_38 ? _GEN_261 : _GEN_229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_301 = _T_38 ? _GEN_262 : _GEN_230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_302 = _T_38 ? _GEN_263 : _GEN_231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_303 = _T_38 ? _GEN_264 : _GEN_232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_304 = _T_38 ? _GEN_265 : _GEN_233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_305 = _T_38 ? _GEN_266 : _GEN_234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_306 = _T_38 ? _GEN_267 : _GEN_235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_307 = _T_38 ? _GEN_268 : _GEN_236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_308 = _T_38 ? _GEN_269 : _GEN_237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_309 = _T_38 ? _GEN_270 : _GEN_238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_310 = _T_38 ? _GEN_271 : _GEN_239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_311 = _T_38 ? _GEN_272 : _GEN_240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_312 = _T_38 ? _GEN_273 : _GEN_241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_313 = _T_38 ? _GEN_274 : _GEN_242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _GEN_314 = _T_38 ? _GEN_275 : _GEN_243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 153:23]
  wire [63:0] _next_reg_T_8 = _GEN_101 & imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:62]
  wire [63:0] _GEN_316 = 5'h1 == rd ? _next_reg_T_8 : _GEN_284; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_317 = 5'h2 == rd ? _next_reg_T_8 : _GEN_285; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_318 = 5'h3 == rd ? _next_reg_T_8 : _GEN_286; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_319 = 5'h4 == rd ? _next_reg_T_8 : _GEN_287; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_320 = 5'h5 == rd ? _next_reg_T_8 : _GEN_288; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_321 = 5'h6 == rd ? _next_reg_T_8 : _GEN_289; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_322 = 5'h7 == rd ? _next_reg_T_8 : _GEN_290; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_323 = 5'h8 == rd ? _next_reg_T_8 : _GEN_291; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_324 = 5'h9 == rd ? _next_reg_T_8 : _GEN_292; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_325 = 5'ha == rd ? _next_reg_T_8 : _GEN_293; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_326 = 5'hb == rd ? _next_reg_T_8 : _GEN_294; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_327 = 5'hc == rd ? _next_reg_T_8 : _GEN_295; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_328 = 5'hd == rd ? _next_reg_T_8 : _GEN_296; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_329 = 5'he == rd ? _next_reg_T_8 : _GEN_297; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_330 = 5'hf == rd ? _next_reg_T_8 : _GEN_298; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_331 = 5'h10 == rd ? _next_reg_T_8 : _GEN_299; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_332 = 5'h11 == rd ? _next_reg_T_8 : _GEN_300; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_333 = 5'h12 == rd ? _next_reg_T_8 : _GEN_301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_334 = 5'h13 == rd ? _next_reg_T_8 : _GEN_302; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_335 = 5'h14 == rd ? _next_reg_T_8 : _GEN_303; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_336 = 5'h15 == rd ? _next_reg_T_8 : _GEN_304; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_337 = 5'h16 == rd ? _next_reg_T_8 : _GEN_305; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_338 = 5'h17 == rd ? _next_reg_T_8 : _GEN_306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_339 = 5'h18 == rd ? _next_reg_T_8 : _GEN_307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_340 = 5'h19 == rd ? _next_reg_T_8 : _GEN_308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_341 = 5'h1a == rd ? _next_reg_T_8 : _GEN_309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_342 = 5'h1b == rd ? _next_reg_T_8 : _GEN_310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_343 = 5'h1c == rd ? _next_reg_T_8 : _GEN_311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_344 = 5'h1d == rd ? _next_reg_T_8 : _GEN_312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_345 = 5'h1e == rd ? _next_reg_T_8 : _GEN_313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_346 = 5'h1f == rd ? _next_reg_T_8 : _GEN_314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:{46,46}]
  wire [63:0] _GEN_355 = _T_44 ? _GEN_316 : _GEN_284; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_356 = _T_44 ? _GEN_317 : _GEN_285; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_357 = _T_44 ? _GEN_318 : _GEN_286; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_358 = _T_44 ? _GEN_319 : _GEN_287; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_359 = _T_44 ? _GEN_320 : _GEN_288; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_360 = _T_44 ? _GEN_321 : _GEN_289; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_361 = _T_44 ? _GEN_322 : _GEN_290; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_362 = _T_44 ? _GEN_323 : _GEN_291; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_363 = _T_44 ? _GEN_324 : _GEN_292; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_364 = _T_44 ? _GEN_325 : _GEN_293; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_365 = _T_44 ? _GEN_326 : _GEN_294; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_366 = _T_44 ? _GEN_327 : _GEN_295; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_367 = _T_44 ? _GEN_328 : _GEN_296; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_368 = _T_44 ? _GEN_329 : _GEN_297; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_369 = _T_44 ? _GEN_330 : _GEN_298; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_370 = _T_44 ? _GEN_331 : _GEN_299; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_371 = _T_44 ? _GEN_332 : _GEN_300; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_372 = _T_44 ? _GEN_333 : _GEN_301; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_373 = _T_44 ? _GEN_334 : _GEN_302; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_374 = _T_44 ? _GEN_335 : _GEN_303; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_375 = _T_44 ? _GEN_336 : _GEN_304; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_376 = _T_44 ? _GEN_337 : _GEN_305; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_377 = _T_44 ? _GEN_338 : _GEN_306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_378 = _T_44 ? _GEN_339 : _GEN_307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_379 = _T_44 ? _GEN_340 : _GEN_308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_380 = _T_44 ? _GEN_341 : _GEN_309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_381 = _T_44 ? _GEN_342 : _GEN_310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_382 = _T_44 ? _GEN_343 : _GEN_311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_383 = _T_44 ? _GEN_344 : _GEN_312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_384 = _T_44 ? _GEN_345 : _GEN_313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _GEN_385 = _T_44 ? _GEN_346 : _GEN_314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 155:22]
  wire [63:0] _next_reg_T_9 = _GEN_101 | imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:62]
  wire [63:0] _GEN_387 = 5'h1 == rd ? _next_reg_T_9 : _GEN_355; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_388 = 5'h2 == rd ? _next_reg_T_9 : _GEN_356; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_389 = 5'h3 == rd ? _next_reg_T_9 : _GEN_357; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_390 = 5'h4 == rd ? _next_reg_T_9 : _GEN_358; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_391 = 5'h5 == rd ? _next_reg_T_9 : _GEN_359; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_392 = 5'h6 == rd ? _next_reg_T_9 : _GEN_360; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_393 = 5'h7 == rd ? _next_reg_T_9 : _GEN_361; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_394 = 5'h8 == rd ? _next_reg_T_9 : _GEN_362; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_395 = 5'h9 == rd ? _next_reg_T_9 : _GEN_363; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_396 = 5'ha == rd ? _next_reg_T_9 : _GEN_364; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_397 = 5'hb == rd ? _next_reg_T_9 : _GEN_365; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_398 = 5'hc == rd ? _next_reg_T_9 : _GEN_366; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_399 = 5'hd == rd ? _next_reg_T_9 : _GEN_367; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_400 = 5'he == rd ? _next_reg_T_9 : _GEN_368; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_401 = 5'hf == rd ? _next_reg_T_9 : _GEN_369; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_402 = 5'h10 == rd ? _next_reg_T_9 : _GEN_370; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_403 = 5'h11 == rd ? _next_reg_T_9 : _GEN_371; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_404 = 5'h12 == rd ? _next_reg_T_9 : _GEN_372; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_405 = 5'h13 == rd ? _next_reg_T_9 : _GEN_373; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_406 = 5'h14 == rd ? _next_reg_T_9 : _GEN_374; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_407 = 5'h15 == rd ? _next_reg_T_9 : _GEN_375; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_408 = 5'h16 == rd ? _next_reg_T_9 : _GEN_376; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_409 = 5'h17 == rd ? _next_reg_T_9 : _GEN_377; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_410 = 5'h18 == rd ? _next_reg_T_9 : _GEN_378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_411 = 5'h19 == rd ? _next_reg_T_9 : _GEN_379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_412 = 5'h1a == rd ? _next_reg_T_9 : _GEN_380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_413 = 5'h1b == rd ? _next_reg_T_9 : _GEN_381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_414 = 5'h1c == rd ? _next_reg_T_9 : _GEN_382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_415 = 5'h1d == rd ? _next_reg_T_9 : _GEN_383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_416 = 5'h1e == rd ? _next_reg_T_9 : _GEN_384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_417 = 5'h1f == rd ? _next_reg_T_9 : _GEN_385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:{46,46}]
  wire [63:0] _GEN_426 = _T_50 ? _GEN_387 : _GEN_355; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_427 = _T_50 ? _GEN_388 : _GEN_356; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_428 = _T_50 ? _GEN_389 : _GEN_357; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_429 = _T_50 ? _GEN_390 : _GEN_358; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_430 = _T_50 ? _GEN_391 : _GEN_359; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_431 = _T_50 ? _GEN_392 : _GEN_360; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_432 = _T_50 ? _GEN_393 : _GEN_361; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_433 = _T_50 ? _GEN_394 : _GEN_362; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_434 = _T_50 ? _GEN_395 : _GEN_363; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_435 = _T_50 ? _GEN_396 : _GEN_364; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_436 = _T_50 ? _GEN_397 : _GEN_365; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_437 = _T_50 ? _GEN_398 : _GEN_366; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_438 = _T_50 ? _GEN_399 : _GEN_367; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_439 = _T_50 ? _GEN_400 : _GEN_368; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_440 = _T_50 ? _GEN_401 : _GEN_369; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_441 = _T_50 ? _GEN_402 : _GEN_370; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_442 = _T_50 ? _GEN_403 : _GEN_371; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_443 = _T_50 ? _GEN_404 : _GEN_372; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_444 = _T_50 ? _GEN_405 : _GEN_373; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_445 = _T_50 ? _GEN_406 : _GEN_374; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_446 = _T_50 ? _GEN_407 : _GEN_375; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_447 = _T_50 ? _GEN_408 : _GEN_376; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_448 = _T_50 ? _GEN_409 : _GEN_377; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_449 = _T_50 ? _GEN_410 : _GEN_378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_450 = _T_50 ? _GEN_411 : _GEN_379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_451 = _T_50 ? _GEN_412 : _GEN_380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_452 = _T_50 ? _GEN_413 : _GEN_381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_453 = _T_50 ? _GEN_414 : _GEN_382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_454 = _T_50 ? _GEN_415 : _GEN_383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_455 = _T_50 ? _GEN_416 : _GEN_384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _GEN_456 = _T_50 ? _GEN_417 : _GEN_385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 156:22]
  wire [63:0] _next_reg_T_10 = _GEN_101 ^ imm; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:62]
  wire [63:0] _GEN_458 = 5'h1 == rd ? _next_reg_T_10 : _GEN_426; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_459 = 5'h2 == rd ? _next_reg_T_10 : _GEN_427; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_460 = 5'h3 == rd ? _next_reg_T_10 : _GEN_428; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_461 = 5'h4 == rd ? _next_reg_T_10 : _GEN_429; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_462 = 5'h5 == rd ? _next_reg_T_10 : _GEN_430; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_463 = 5'h6 == rd ? _next_reg_T_10 : _GEN_431; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_464 = 5'h7 == rd ? _next_reg_T_10 : _GEN_432; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_465 = 5'h8 == rd ? _next_reg_T_10 : _GEN_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_466 = 5'h9 == rd ? _next_reg_T_10 : _GEN_434; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_467 = 5'ha == rd ? _next_reg_T_10 : _GEN_435; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_468 = 5'hb == rd ? _next_reg_T_10 : _GEN_436; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_469 = 5'hc == rd ? _next_reg_T_10 : _GEN_437; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_470 = 5'hd == rd ? _next_reg_T_10 : _GEN_438; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_471 = 5'he == rd ? _next_reg_T_10 : _GEN_439; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_472 = 5'hf == rd ? _next_reg_T_10 : _GEN_440; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_473 = 5'h10 == rd ? _next_reg_T_10 : _GEN_441; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_474 = 5'h11 == rd ? _next_reg_T_10 : _GEN_442; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_475 = 5'h12 == rd ? _next_reg_T_10 : _GEN_443; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_476 = 5'h13 == rd ? _next_reg_T_10 : _GEN_444; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_477 = 5'h14 == rd ? _next_reg_T_10 : _GEN_445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_478 = 5'h15 == rd ? _next_reg_T_10 : _GEN_446; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_479 = 5'h16 == rd ? _next_reg_T_10 : _GEN_447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_480 = 5'h17 == rd ? _next_reg_T_10 : _GEN_448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_481 = 5'h18 == rd ? _next_reg_T_10 : _GEN_449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_482 = 5'h19 == rd ? _next_reg_T_10 : _GEN_450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_483 = 5'h1a == rd ? _next_reg_T_10 : _GEN_451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_484 = 5'h1b == rd ? _next_reg_T_10 : _GEN_452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_485 = 5'h1c == rd ? _next_reg_T_10 : _GEN_453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_486 = 5'h1d == rd ? _next_reg_T_10 : _GEN_454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_487 = 5'h1e == rd ? _next_reg_T_10 : _GEN_455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_488 = 5'h1f == rd ? _next_reg_T_10 : _GEN_456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:{46,46}]
  wire [63:0] _GEN_497 = _T_56 ? _GEN_458 : _GEN_426; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_498 = _T_56 ? _GEN_459 : _GEN_427; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_499 = _T_56 ? _GEN_460 : _GEN_428; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_500 = _T_56 ? _GEN_461 : _GEN_429; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_501 = _T_56 ? _GEN_462 : _GEN_430; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_502 = _T_56 ? _GEN_463 : _GEN_431; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_503 = _T_56 ? _GEN_464 : _GEN_432; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_504 = _T_56 ? _GEN_465 : _GEN_433; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_505 = _T_56 ? _GEN_466 : _GEN_434; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_506 = _T_56 ? _GEN_467 : _GEN_435; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_507 = _T_56 ? _GEN_468 : _GEN_436; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_508 = _T_56 ? _GEN_469 : _GEN_437; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_509 = _T_56 ? _GEN_470 : _GEN_438; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_510 = _T_56 ? _GEN_471 : _GEN_439; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_511 = _T_56 ? _GEN_472 : _GEN_440; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_512 = _T_56 ? _GEN_473 : _GEN_441; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_513 = _T_56 ? _GEN_474 : _GEN_442; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_514 = _T_56 ? _GEN_475 : _GEN_443; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_515 = _T_56 ? _GEN_476 : _GEN_444; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_516 = _T_56 ? _GEN_477 : _GEN_445; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_517 = _T_56 ? _GEN_478 : _GEN_446; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_518 = _T_56 ? _GEN_479 : _GEN_447; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_519 = _T_56 ? _GEN_480 : _GEN_448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_520 = _T_56 ? _GEN_481 : _GEN_449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_521 = _T_56 ? _GEN_482 : _GEN_450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_522 = _T_56 ? _GEN_483 : _GEN_451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_523 = _T_56 ? _GEN_484 : _GEN_452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_524 = _T_56 ? _GEN_485 : _GEN_453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_525 = _T_56 ? _GEN_486 : _GEN_454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_526 = _T_56 ? _GEN_487 : _GEN_455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [63:0] _GEN_527 = _T_56 ? _GEN_488 : _GEN_456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 157:22]
  wire [94:0] _GEN_0 = {{31'd0}, _GEN_101}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:62]
  wire [94:0] _next_reg_T_12 = _GEN_0 << imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:62]
  wire [63:0] _GEN_529 = 5'h1 == rd ? _next_reg_T_12[63:0] : _GEN_497; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_530 = 5'h2 == rd ? _next_reg_T_12[63:0] : _GEN_498; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_531 = 5'h3 == rd ? _next_reg_T_12[63:0] : _GEN_499; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_532 = 5'h4 == rd ? _next_reg_T_12[63:0] : _GEN_500; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_533 = 5'h5 == rd ? _next_reg_T_12[63:0] : _GEN_501; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_534 = 5'h6 == rd ? _next_reg_T_12[63:0] : _GEN_502; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_535 = 5'h7 == rd ? _next_reg_T_12[63:0] : _GEN_503; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_536 = 5'h8 == rd ? _next_reg_T_12[63:0] : _GEN_504; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_537 = 5'h9 == rd ? _next_reg_T_12[63:0] : _GEN_505; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_538 = 5'ha == rd ? _next_reg_T_12[63:0] : _GEN_506; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_539 = 5'hb == rd ? _next_reg_T_12[63:0] : _GEN_507; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_540 = 5'hc == rd ? _next_reg_T_12[63:0] : _GEN_508; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_541 = 5'hd == rd ? _next_reg_T_12[63:0] : _GEN_509; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_542 = 5'he == rd ? _next_reg_T_12[63:0] : _GEN_510; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_543 = 5'hf == rd ? _next_reg_T_12[63:0] : _GEN_511; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_544 = 5'h10 == rd ? _next_reg_T_12[63:0] : _GEN_512; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_545 = 5'h11 == rd ? _next_reg_T_12[63:0] : _GEN_513; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_546 = 5'h12 == rd ? _next_reg_T_12[63:0] : _GEN_514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_547 = 5'h13 == rd ? _next_reg_T_12[63:0] : _GEN_515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_548 = 5'h14 == rd ? _next_reg_T_12[63:0] : _GEN_516; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_549 = 5'h15 == rd ? _next_reg_T_12[63:0] : _GEN_517; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_550 = 5'h16 == rd ? _next_reg_T_12[63:0] : _GEN_518; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_551 = 5'h17 == rd ? _next_reg_T_12[63:0] : _GEN_519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_552 = 5'h18 == rd ? _next_reg_T_12[63:0] : _GEN_520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_553 = 5'h19 == rd ? _next_reg_T_12[63:0] : _GEN_521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_554 = 5'h1a == rd ? _next_reg_T_12[63:0] : _GEN_522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_555 = 5'h1b == rd ? _next_reg_T_12[63:0] : _GEN_523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_556 = 5'h1c == rd ? _next_reg_T_12[63:0] : _GEN_524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_557 = 5'h1d == rd ? _next_reg_T_12[63:0] : _GEN_525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_558 = 5'h1e == rd ? _next_reg_T_12[63:0] : _GEN_526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_559 = 5'h1f == rd ? _next_reg_T_12[63:0] : _GEN_527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:{46,46}]
  wire [63:0] _GEN_568 = _T_726 ? _GEN_529 : _GEN_497; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_569 = _T_726 ? _GEN_530 : _GEN_498; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_570 = _T_726 ? _GEN_531 : _GEN_499; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_571 = _T_726 ? _GEN_532 : _GEN_500; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_572 = _T_726 ? _GEN_533 : _GEN_501; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_573 = _T_726 ? _GEN_534 : _GEN_502; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_574 = _T_726 ? _GEN_535 : _GEN_503; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_575 = _T_726 ? _GEN_536 : _GEN_504; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_576 = _T_726 ? _GEN_537 : _GEN_505; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_577 = _T_726 ? _GEN_538 : _GEN_506; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_578 = _T_726 ? _GEN_539 : _GEN_507; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_579 = _T_726 ? _GEN_540 : _GEN_508; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_580 = _T_726 ? _GEN_541 : _GEN_509; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_581 = _T_726 ? _GEN_542 : _GEN_510; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_582 = _T_726 ? _GEN_543 : _GEN_511; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_583 = _T_726 ? _GEN_544 : _GEN_512; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_584 = _T_726 ? _GEN_545 : _GEN_513; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_585 = _T_726 ? _GEN_546 : _GEN_514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_586 = _T_726 ? _GEN_547 : _GEN_515; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_587 = _T_726 ? _GEN_548 : _GEN_516; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_588 = _T_726 ? _GEN_549 : _GEN_517; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_589 = _T_726 ? _GEN_550 : _GEN_518; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_590 = _T_726 ? _GEN_551 : _GEN_519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_591 = _T_726 ? _GEN_552 : _GEN_520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_592 = _T_726 ? _GEN_553 : _GEN_521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_593 = _T_726 ? _GEN_554 : _GEN_522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_594 = _T_726 ? _GEN_555 : _GEN_523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_595 = _T_726 ? _GEN_556 : _GEN_524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_596 = _T_726 ? _GEN_557 : _GEN_525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_597 = _T_726 ? _GEN_558 : _GEN_526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _GEN_598 = _T_726 ? _GEN_559 : _GEN_527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 159:22]
  wire [63:0] _next_reg_T_14 = _GEN_101 >> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:62]
  wire [63:0] _GEN_600 = 5'h1 == rd ? _next_reg_T_14 : _GEN_568; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_601 = 5'h2 == rd ? _next_reg_T_14 : _GEN_569; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_602 = 5'h3 == rd ? _next_reg_T_14 : _GEN_570; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_603 = 5'h4 == rd ? _next_reg_T_14 : _GEN_571; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_604 = 5'h5 == rd ? _next_reg_T_14 : _GEN_572; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_605 = 5'h6 == rd ? _next_reg_T_14 : _GEN_573; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_606 = 5'h7 == rd ? _next_reg_T_14 : _GEN_574; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_607 = 5'h8 == rd ? _next_reg_T_14 : _GEN_575; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_608 = 5'h9 == rd ? _next_reg_T_14 : _GEN_576; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_609 = 5'ha == rd ? _next_reg_T_14 : _GEN_577; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_610 = 5'hb == rd ? _next_reg_T_14 : _GEN_578; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_611 = 5'hc == rd ? _next_reg_T_14 : _GEN_579; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_612 = 5'hd == rd ? _next_reg_T_14 : _GEN_580; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_613 = 5'he == rd ? _next_reg_T_14 : _GEN_581; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_614 = 5'hf == rd ? _next_reg_T_14 : _GEN_582; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_615 = 5'h10 == rd ? _next_reg_T_14 : _GEN_583; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_616 = 5'h11 == rd ? _next_reg_T_14 : _GEN_584; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_617 = 5'h12 == rd ? _next_reg_T_14 : _GEN_585; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_618 = 5'h13 == rd ? _next_reg_T_14 : _GEN_586; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_619 = 5'h14 == rd ? _next_reg_T_14 : _GEN_587; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_620 = 5'h15 == rd ? _next_reg_T_14 : _GEN_588; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_621 = 5'h16 == rd ? _next_reg_T_14 : _GEN_589; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_622 = 5'h17 == rd ? _next_reg_T_14 : _GEN_590; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_623 = 5'h18 == rd ? _next_reg_T_14 : _GEN_591; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_624 = 5'h19 == rd ? _next_reg_T_14 : _GEN_592; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_625 = 5'h1a == rd ? _next_reg_T_14 : _GEN_593; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_626 = 5'h1b == rd ? _next_reg_T_14 : _GEN_594; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_627 = 5'h1c == rd ? _next_reg_T_14 : _GEN_595; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_628 = 5'h1d == rd ? _next_reg_T_14 : _GEN_596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_629 = 5'h1e == rd ? _next_reg_T_14 : _GEN_597; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_630 = 5'h1f == rd ? _next_reg_T_14 : _GEN_598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:{46,46}]
  wire [63:0] _GEN_639 = _T_732 ? _GEN_600 : _GEN_568; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_640 = _T_732 ? _GEN_601 : _GEN_569; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_641 = _T_732 ? _GEN_602 : _GEN_570; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_642 = _T_732 ? _GEN_603 : _GEN_571; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_643 = _T_732 ? _GEN_604 : _GEN_572; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_644 = _T_732 ? _GEN_605 : _GEN_573; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_645 = _T_732 ? _GEN_606 : _GEN_574; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_646 = _T_732 ? _GEN_607 : _GEN_575; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_647 = _T_732 ? _GEN_608 : _GEN_576; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_648 = _T_732 ? _GEN_609 : _GEN_577; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_649 = _T_732 ? _GEN_610 : _GEN_578; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_650 = _T_732 ? _GEN_611 : _GEN_579; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_651 = _T_732 ? _GEN_612 : _GEN_580; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_652 = _T_732 ? _GEN_613 : _GEN_581; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_653 = _T_732 ? _GEN_614 : _GEN_582; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_654 = _T_732 ? _GEN_615 : _GEN_583; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_655 = _T_732 ? _GEN_616 : _GEN_584; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_656 = _T_732 ? _GEN_617 : _GEN_585; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_657 = _T_732 ? _GEN_618 : _GEN_586; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_658 = _T_732 ? _GEN_619 : _GEN_587; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_659 = _T_732 ? _GEN_620 : _GEN_588; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_660 = _T_732 ? _GEN_621 : _GEN_589; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_661 = _T_732 ? _GEN_622 : _GEN_590; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_662 = _T_732 ? _GEN_623 : _GEN_591; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_663 = _T_732 ? _GEN_624 : _GEN_592; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_664 = _T_732 ? _GEN_625 : _GEN_593; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_665 = _T_732 ? _GEN_626 : _GEN_594; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_666 = _T_732 ? _GEN_627 : _GEN_595; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_667 = _T_732 ? _GEN_628 : _GEN_596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_668 = _T_732 ? _GEN_629 : _GEN_597; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _GEN_669 = _T_732 ? _GEN_630 : _GEN_598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 160:22]
  wire [63:0] _next_reg_T_18 = $signed(_T_325) >>> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:84]
  wire [63:0] _GEN_671 = 5'h1 == rd ? _next_reg_T_18 : _GEN_639; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_672 = 5'h2 == rd ? _next_reg_T_18 : _GEN_640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_673 = 5'h3 == rd ? _next_reg_T_18 : _GEN_641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_674 = 5'h4 == rd ? _next_reg_T_18 : _GEN_642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_675 = 5'h5 == rd ? _next_reg_T_18 : _GEN_643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_676 = 5'h6 == rd ? _next_reg_T_18 : _GEN_644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_677 = 5'h7 == rd ? _next_reg_T_18 : _GEN_645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_678 = 5'h8 == rd ? _next_reg_T_18 : _GEN_646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_679 = 5'h9 == rd ? _next_reg_T_18 : _GEN_647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_680 = 5'ha == rd ? _next_reg_T_18 : _GEN_648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_681 = 5'hb == rd ? _next_reg_T_18 : _GEN_649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_682 = 5'hc == rd ? _next_reg_T_18 : _GEN_650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_683 = 5'hd == rd ? _next_reg_T_18 : _GEN_651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_684 = 5'he == rd ? _next_reg_T_18 : _GEN_652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_685 = 5'hf == rd ? _next_reg_T_18 : _GEN_653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_686 = 5'h10 == rd ? _next_reg_T_18 : _GEN_654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_687 = 5'h11 == rd ? _next_reg_T_18 : _GEN_655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_688 = 5'h12 == rd ? _next_reg_T_18 : _GEN_656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_689 = 5'h13 == rd ? _next_reg_T_18 : _GEN_657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_690 = 5'h14 == rd ? _next_reg_T_18 : _GEN_658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_691 = 5'h15 == rd ? _next_reg_T_18 : _GEN_659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_692 = 5'h16 == rd ? _next_reg_T_18 : _GEN_660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_693 = 5'h17 == rd ? _next_reg_T_18 : _GEN_661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_694 = 5'h18 == rd ? _next_reg_T_18 : _GEN_662; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_695 = 5'h19 == rd ? _next_reg_T_18 : _GEN_663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_696 = 5'h1a == rd ? _next_reg_T_18 : _GEN_664; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_697 = 5'h1b == rd ? _next_reg_T_18 : _GEN_665; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_698 = 5'h1c == rd ? _next_reg_T_18 : _GEN_666; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_699 = 5'h1d == rd ? _next_reg_T_18 : _GEN_667; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_700 = 5'h1e == rd ? _next_reg_T_18 : _GEN_668; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_701 = 5'h1f == rd ? _next_reg_T_18 : _GEN_669; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:{46,46}]
  wire [63:0] _GEN_710 = _T_738 ? _GEN_671 : _GEN_639; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_711 = _T_738 ? _GEN_672 : _GEN_640; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_712 = _T_738 ? _GEN_673 : _GEN_641; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_713 = _T_738 ? _GEN_674 : _GEN_642; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_714 = _T_738 ? _GEN_675 : _GEN_643; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_715 = _T_738 ? _GEN_676 : _GEN_644; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_716 = _T_738 ? _GEN_677 : _GEN_645; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_717 = _T_738 ? _GEN_678 : _GEN_646; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_718 = _T_738 ? _GEN_679 : _GEN_647; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_719 = _T_738 ? _GEN_680 : _GEN_648; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_720 = _T_738 ? _GEN_681 : _GEN_649; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_721 = _T_738 ? _GEN_682 : _GEN_650; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_722 = _T_738 ? _GEN_683 : _GEN_651; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_723 = _T_738 ? _GEN_684 : _GEN_652; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_724 = _T_738 ? _GEN_685 : _GEN_653; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_725 = _T_738 ? _GEN_686 : _GEN_654; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_726 = _T_738 ? _GEN_687 : _GEN_655; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_727 = _T_738 ? _GEN_688 : _GEN_656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_728 = _T_738 ? _GEN_689 : _GEN_657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_729 = _T_738 ? _GEN_690 : _GEN_658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_730 = _T_738 ? _GEN_691 : _GEN_659; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_731 = _T_738 ? _GEN_692 : _GEN_660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_732 = _T_738 ? _GEN_693 : _GEN_661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_733 = _T_738 ? _GEN_694 : _GEN_662; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_734 = _T_738 ? _GEN_695 : _GEN_663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_735 = _T_738 ? _GEN_696 : _GEN_664; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_736 = _T_738 ? _GEN_697 : _GEN_665; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_737 = _T_738 ? _GEN_698 : _GEN_666; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_738 = _T_738 ? _GEN_699 : _GEN_667; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_739 = _T_738 ? _GEN_700 : _GEN_668; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_740 = _T_738 ? _GEN_701 : _GEN_669; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 161:22]
  wire [63:0] _GEN_742 = 5'h1 == rd ? imm : _GEN_710; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_743 = 5'h2 == rd ? imm : _GEN_711; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_744 = 5'h3 == rd ? imm : _GEN_712; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_745 = 5'h4 == rd ? imm : _GEN_713; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_746 = 5'h5 == rd ? imm : _GEN_714; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_747 = 5'h6 == rd ? imm : _GEN_715; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_748 = 5'h7 == rd ? imm : _GEN_716; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_749 = 5'h8 == rd ? imm : _GEN_717; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_750 = 5'h9 == rd ? imm : _GEN_718; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_751 = 5'ha == rd ? imm : _GEN_719; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_752 = 5'hb == rd ? imm : _GEN_720; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_753 = 5'hc == rd ? imm : _GEN_721; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_754 = 5'hd == rd ? imm : _GEN_722; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_755 = 5'he == rd ? imm : _GEN_723; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_756 = 5'hf == rd ? imm : _GEN_724; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_757 = 5'h10 == rd ? imm : _GEN_725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_758 = 5'h11 == rd ? imm : _GEN_726; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_759 = 5'h12 == rd ? imm : _GEN_727; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_760 = 5'h13 == rd ? imm : _GEN_728; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_761 = 5'h14 == rd ? imm : _GEN_729; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_762 = 5'h15 == rd ? imm : _GEN_730; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_763 = 5'h16 == rd ? imm : _GEN_731; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_764 = 5'h17 == rd ? imm : _GEN_732; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_765 = 5'h18 == rd ? imm : _GEN_733; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_766 = 5'h19 == rd ? imm : _GEN_734; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_767 = 5'h1a == rd ? imm : _GEN_735; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_768 = 5'h1b == rd ? imm : _GEN_736; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_769 = 5'h1c == rd ? imm : _GEN_737; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_770 = 5'h1d == rd ? imm : _GEN_738; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_771 = 5'h1e == rd ? imm : _GEN_739; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_772 = 5'h1f == rd ? imm : _GEN_740; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:{45,45}]
  wire [63:0] _GEN_779 = _T_80 ? _GEN_742 : _GEN_710; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_780 = _T_80 ? _GEN_743 : _GEN_711; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_781 = _T_80 ? _GEN_744 : _GEN_712; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_782 = _T_80 ? _GEN_745 : _GEN_713; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_783 = _T_80 ? _GEN_746 : _GEN_714; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_784 = _T_80 ? _GEN_747 : _GEN_715; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_785 = _T_80 ? _GEN_748 : _GEN_716; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_786 = _T_80 ? _GEN_749 : _GEN_717; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_787 = _T_80 ? _GEN_750 : _GEN_718; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_788 = _T_80 ? _GEN_751 : _GEN_719; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_789 = _T_80 ? _GEN_752 : _GEN_720; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_790 = _T_80 ? _GEN_753 : _GEN_721; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_791 = _T_80 ? _GEN_754 : _GEN_722; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_792 = _T_80 ? _GEN_755 : _GEN_723; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_793 = _T_80 ? _GEN_756 : _GEN_724; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_794 = _T_80 ? _GEN_757 : _GEN_725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_795 = _T_80 ? _GEN_758 : _GEN_726; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_796 = _T_80 ? _GEN_759 : _GEN_727; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_797 = _T_80 ? _GEN_760 : _GEN_728; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_798 = _T_80 ? _GEN_761 : _GEN_729; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_799 = _T_80 ? _GEN_762 : _GEN_730; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_800 = _T_80 ? _GEN_763 : _GEN_731; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_801 = _T_80 ? _GEN_764 : _GEN_732; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_802 = _T_80 ? _GEN_765 : _GEN_733; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_803 = _T_80 ? _GEN_766 : _GEN_734; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_804 = _T_80 ? _GEN_767 : _GEN_735; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_805 = _T_80 ? _GEN_768 : _GEN_736; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_806 = _T_80 ? _GEN_769 : _GEN_737; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_807 = _T_80 ? _GEN_770 : _GEN_738; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_808 = _T_80 ? _GEN_771 : _GEN_739; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_809 = _T_80 ? _GEN_772 : _GEN_740; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 163:21]
  wire [63:0] _GEN_811 = 5'h1 == rd ? _T_359 : _GEN_779; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_812 = 5'h2 == rd ? _T_359 : _GEN_780; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_813 = 5'h3 == rd ? _T_359 : _GEN_781; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_814 = 5'h4 == rd ? _T_359 : _GEN_782; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_815 = 5'h5 == rd ? _T_359 : _GEN_783; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_816 = 5'h6 == rd ? _T_359 : _GEN_784; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_817 = 5'h7 == rd ? _T_359 : _GEN_785; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_818 = 5'h8 == rd ? _T_359 : _GEN_786; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_819 = 5'h9 == rd ? _T_359 : _GEN_787; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_820 = 5'ha == rd ? _T_359 : _GEN_788; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_821 = 5'hb == rd ? _T_359 : _GEN_789; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_822 = 5'hc == rd ? _T_359 : _GEN_790; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_823 = 5'hd == rd ? _T_359 : _GEN_791; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_824 = 5'he == rd ? _T_359 : _GEN_792; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_825 = 5'hf == rd ? _T_359 : _GEN_793; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_826 = 5'h10 == rd ? _T_359 : _GEN_794; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_827 = 5'h11 == rd ? _T_359 : _GEN_795; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_828 = 5'h12 == rd ? _T_359 : _GEN_796; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_829 = 5'h13 == rd ? _T_359 : _GEN_797; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_830 = 5'h14 == rd ? _T_359 : _GEN_798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_831 = 5'h15 == rd ? _T_359 : _GEN_799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_832 = 5'h16 == rd ? _T_359 : _GEN_800; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_833 = 5'h17 == rd ? _T_359 : _GEN_801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_834 = 5'h18 == rd ? _T_359 : _GEN_802; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_835 = 5'h19 == rd ? _T_359 : _GEN_803; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_836 = 5'h1a == rd ? _T_359 : _GEN_804; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_837 = 5'h1b == rd ? _T_359 : _GEN_805; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_838 = 5'h1c == rd ? _T_359 : _GEN_806; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_839 = 5'h1d == rd ? _T_359 : _GEN_807; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_840 = 5'h1e == rd ? _T_359 : _GEN_808; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_841 = 5'h1f == rd ? _T_359 : _GEN_809; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:{47,47}]
  wire [63:0] _GEN_848 = _T_84 ? _GEN_811 : _GEN_779; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_849 = _T_84 ? _GEN_812 : _GEN_780; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_850 = _T_84 ? _GEN_813 : _GEN_781; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_851 = _T_84 ? _GEN_814 : _GEN_782; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_852 = _T_84 ? _GEN_815 : _GEN_783; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_853 = _T_84 ? _GEN_816 : _GEN_784; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_854 = _T_84 ? _GEN_817 : _GEN_785; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_855 = _T_84 ? _GEN_818 : _GEN_786; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_856 = _T_84 ? _GEN_819 : _GEN_787; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_857 = _T_84 ? _GEN_820 : _GEN_788; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_858 = _T_84 ? _GEN_821 : _GEN_789; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_859 = _T_84 ? _GEN_822 : _GEN_790; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_860 = _T_84 ? _GEN_823 : _GEN_791; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_861 = _T_84 ? _GEN_824 : _GEN_792; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_862 = _T_84 ? _GEN_825 : _GEN_793; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_863 = _T_84 ? _GEN_826 : _GEN_794; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_864 = _T_84 ? _GEN_827 : _GEN_795; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_865 = _T_84 ? _GEN_828 : _GEN_796; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_866 = _T_84 ? _GEN_829 : _GEN_797; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_867 = _T_84 ? _GEN_830 : _GEN_798; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_868 = _T_84 ? _GEN_831 : _GEN_799; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_869 = _T_84 ? _GEN_832 : _GEN_800; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_870 = _T_84 ? _GEN_833 : _GEN_801; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_871 = _T_84 ? _GEN_834 : _GEN_802; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_872 = _T_84 ? _GEN_835 : _GEN_803; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_873 = _T_84 ? _GEN_836 : _GEN_804; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_874 = _T_84 ? _GEN_837 : _GEN_805; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_875 = _T_84 ? _GEN_838 : _GEN_806; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_876 = _T_84 ? _GEN_839 : _GEN_807; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_877 = _T_84 ? _GEN_840 : _GEN_808; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _GEN_878 = _T_84 ? _GEN_841 : _GEN_809; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 165:23]
  wire [63:0] _next_reg_T_22 = _GEN_101 + _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:62]
  wire [63:0] _GEN_912 = 5'h1 == rd ? _next_reg_T_22 : _GEN_848; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_913 = 5'h2 == rd ? _next_reg_T_22 : _GEN_849; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_914 = 5'h3 == rd ? _next_reg_T_22 : _GEN_850; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_915 = 5'h4 == rd ? _next_reg_T_22 : _GEN_851; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_916 = 5'h5 == rd ? _next_reg_T_22 : _GEN_852; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_917 = 5'h6 == rd ? _next_reg_T_22 : _GEN_853; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_918 = 5'h7 == rd ? _next_reg_T_22 : _GEN_854; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_919 = 5'h8 == rd ? _next_reg_T_22 : _GEN_855; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_920 = 5'h9 == rd ? _next_reg_T_22 : _GEN_856; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_921 = 5'ha == rd ? _next_reg_T_22 : _GEN_857; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_922 = 5'hb == rd ? _next_reg_T_22 : _GEN_858; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_923 = 5'hc == rd ? _next_reg_T_22 : _GEN_859; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_924 = 5'hd == rd ? _next_reg_T_22 : _GEN_860; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_925 = 5'he == rd ? _next_reg_T_22 : _GEN_861; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_926 = 5'hf == rd ? _next_reg_T_22 : _GEN_862; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_927 = 5'h10 == rd ? _next_reg_T_22 : _GEN_863; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_928 = 5'h11 == rd ? _next_reg_T_22 : _GEN_864; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_929 = 5'h12 == rd ? _next_reg_T_22 : _GEN_865; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_930 = 5'h13 == rd ? _next_reg_T_22 : _GEN_866; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_931 = 5'h14 == rd ? _next_reg_T_22 : _GEN_867; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_932 = 5'h15 == rd ? _next_reg_T_22 : _GEN_868; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_933 = 5'h16 == rd ? _next_reg_T_22 : _GEN_869; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_934 = 5'h17 == rd ? _next_reg_T_22 : _GEN_870; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_935 = 5'h18 == rd ? _next_reg_T_22 : _GEN_871; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_936 = 5'h19 == rd ? _next_reg_T_22 : _GEN_872; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_937 = 5'h1a == rd ? _next_reg_T_22 : _GEN_873; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_938 = 5'h1b == rd ? _next_reg_T_22 : _GEN_874; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_939 = 5'h1c == rd ? _next_reg_T_22 : _GEN_875; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_940 = 5'h1d == rd ? _next_reg_T_22 : _GEN_876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_941 = 5'h1e == rd ? _next_reg_T_22 : _GEN_877; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_942 = 5'h1f == rd ? _next_reg_T_22 : _GEN_878; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:{46,46}]
  wire [63:0] _GEN_951 = _T_88 ? _GEN_912 : _GEN_848; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_952 = _T_88 ? _GEN_913 : _GEN_849; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_953 = _T_88 ? _GEN_914 : _GEN_850; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_954 = _T_88 ? _GEN_915 : _GEN_851; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_955 = _T_88 ? _GEN_916 : _GEN_852; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_956 = _T_88 ? _GEN_917 : _GEN_853; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_957 = _T_88 ? _GEN_918 : _GEN_854; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_958 = _T_88 ? _GEN_919 : _GEN_855; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_959 = _T_88 ? _GEN_920 : _GEN_856; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_960 = _T_88 ? _GEN_921 : _GEN_857; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_961 = _T_88 ? _GEN_922 : _GEN_858; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_962 = _T_88 ? _GEN_923 : _GEN_859; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_963 = _T_88 ? _GEN_924 : _GEN_860; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_964 = _T_88 ? _GEN_925 : _GEN_861; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_965 = _T_88 ? _GEN_926 : _GEN_862; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_966 = _T_88 ? _GEN_927 : _GEN_863; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_967 = _T_88 ? _GEN_928 : _GEN_864; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_968 = _T_88 ? _GEN_929 : _GEN_865; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_969 = _T_88 ? _GEN_930 : _GEN_866; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_970 = _T_88 ? _GEN_931 : _GEN_867; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_971 = _T_88 ? _GEN_932 : _GEN_868; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_972 = _T_88 ? _GEN_933 : _GEN_869; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_973 = _T_88 ? _GEN_934 : _GEN_870; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_974 = _T_88 ? _GEN_935 : _GEN_871; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_975 = _T_88 ? _GEN_936 : _GEN_872; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_976 = _T_88 ? _GEN_937 : _GEN_873; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_977 = _T_88 ? _GEN_938 : _GEN_874; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_978 = _T_88 ? _GEN_939 : _GEN_875; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_979 = _T_88 ? _GEN_940 : _GEN_876; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_980 = _T_88 ? _GEN_941 : _GEN_877; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _GEN_981 = _T_88 ? _GEN_942 : _GEN_878; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 168:22]
  wire [63:0] _next_reg_rd_11 = {{63'd0}, _T_271}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_983 = 5'h1 == rd ? _next_reg_rd_11 : _GEN_951; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_984 = 5'h2 == rd ? _next_reg_rd_11 : _GEN_952; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_985 = 5'h3 == rd ? _next_reg_rd_11 : _GEN_953; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_986 = 5'h4 == rd ? _next_reg_rd_11 : _GEN_954; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_987 = 5'h5 == rd ? _next_reg_rd_11 : _GEN_955; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_988 = 5'h6 == rd ? _next_reg_rd_11 : _GEN_956; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_989 = 5'h7 == rd ? _next_reg_rd_11 : _GEN_957; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_990 = 5'h8 == rd ? _next_reg_rd_11 : _GEN_958; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_991 = 5'h9 == rd ? _next_reg_rd_11 : _GEN_959; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_992 = 5'ha == rd ? _next_reg_rd_11 : _GEN_960; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_993 = 5'hb == rd ? _next_reg_rd_11 : _GEN_961; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_994 = 5'hc == rd ? _next_reg_rd_11 : _GEN_962; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_995 = 5'hd == rd ? _next_reg_rd_11 : _GEN_963; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_996 = 5'he == rd ? _next_reg_rd_11 : _GEN_964; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_997 = 5'hf == rd ? _next_reg_rd_11 : _GEN_965; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_998 = 5'h10 == rd ? _next_reg_rd_11 : _GEN_966; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_999 = 5'h11 == rd ? _next_reg_rd_11 : _GEN_967; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_1000 = 5'h12 == rd ? _next_reg_rd_11 : _GEN_968; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_1001 = 5'h13 == rd ? _next_reg_rd_11 : _GEN_969; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_1002 = 5'h14 == rd ? _next_reg_rd_11 : _GEN_970; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_1003 = 5'h15 == rd ? _next_reg_rd_11 : _GEN_971; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_1004 = 5'h16 == rd ? _next_reg_rd_11 : _GEN_972; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_1005 = 5'h17 == rd ? _next_reg_rd_11 : _GEN_973; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_1006 = 5'h18 == rd ? _next_reg_rd_11 : _GEN_974; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_1007 = 5'h19 == rd ? _next_reg_rd_11 : _GEN_975; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_1008 = 5'h1a == rd ? _next_reg_rd_11 : _GEN_976; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_1009 = 5'h1b == rd ? _next_reg_rd_11 : _GEN_977; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_1010 = 5'h1c == rd ? _next_reg_rd_11 : _GEN_978; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_1011 = 5'h1d == rd ? _next_reg_rd_11 : _GEN_979; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_1012 = 5'h1e == rd ? _next_reg_rd_11 : _GEN_980; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_1013 = 5'h1f == rd ? _next_reg_rd_11 : _GEN_981; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:{46,46}]
  wire [63:0] _GEN_1022 = _T_95 ? _GEN_983 : _GEN_951; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1023 = _T_95 ? _GEN_984 : _GEN_952; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1024 = _T_95 ? _GEN_985 : _GEN_953; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1025 = _T_95 ? _GEN_986 : _GEN_954; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1026 = _T_95 ? _GEN_987 : _GEN_955; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1027 = _T_95 ? _GEN_988 : _GEN_956; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1028 = _T_95 ? _GEN_989 : _GEN_957; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1029 = _T_95 ? _GEN_990 : _GEN_958; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1030 = _T_95 ? _GEN_991 : _GEN_959; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1031 = _T_95 ? _GEN_992 : _GEN_960; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1032 = _T_95 ? _GEN_993 : _GEN_961; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1033 = _T_95 ? _GEN_994 : _GEN_962; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1034 = _T_95 ? _GEN_995 : _GEN_963; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1035 = _T_95 ? _GEN_996 : _GEN_964; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1036 = _T_95 ? _GEN_997 : _GEN_965; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1037 = _T_95 ? _GEN_998 : _GEN_966; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1038 = _T_95 ? _GEN_999 : _GEN_967; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1039 = _T_95 ? _GEN_1000 : _GEN_968; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1040 = _T_95 ? _GEN_1001 : _GEN_969; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1041 = _T_95 ? _GEN_1002 : _GEN_970; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1042 = _T_95 ? _GEN_1003 : _GEN_971; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1043 = _T_95 ? _GEN_1004 : _GEN_972; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1044 = _T_95 ? _GEN_1005 : _GEN_973; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1045 = _T_95 ? _GEN_1006 : _GEN_974; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1046 = _T_95 ? _GEN_1007 : _GEN_975; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1047 = _T_95 ? _GEN_1008 : _GEN_976; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1048 = _T_95 ? _GEN_1009 : _GEN_977; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1049 = _T_95 ? _GEN_1010 : _GEN_978; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1050 = _T_95 ? _GEN_1011 : _GEN_979; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1051 = _T_95 ? _GEN_1012 : _GEN_980; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _GEN_1052 = _T_95 ? _GEN_1013 : _GEN_981; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 169:22]
  wire [63:0] _next_reg_rd_12 = {{63'd0}, _T_298}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1054 = 5'h1 == rd ? _next_reg_rd_12 : _GEN_1022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1055 = 5'h2 == rd ? _next_reg_rd_12 : _GEN_1023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1056 = 5'h3 == rd ? _next_reg_rd_12 : _GEN_1024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1057 = 5'h4 == rd ? _next_reg_rd_12 : _GEN_1025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1058 = 5'h5 == rd ? _next_reg_rd_12 : _GEN_1026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1059 = 5'h6 == rd ? _next_reg_rd_12 : _GEN_1027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1060 = 5'h7 == rd ? _next_reg_rd_12 : _GEN_1028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1061 = 5'h8 == rd ? _next_reg_rd_12 : _GEN_1029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1062 = 5'h9 == rd ? _next_reg_rd_12 : _GEN_1030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1063 = 5'ha == rd ? _next_reg_rd_12 : _GEN_1031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1064 = 5'hb == rd ? _next_reg_rd_12 : _GEN_1032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1065 = 5'hc == rd ? _next_reg_rd_12 : _GEN_1033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1066 = 5'hd == rd ? _next_reg_rd_12 : _GEN_1034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1067 = 5'he == rd ? _next_reg_rd_12 : _GEN_1035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1068 = 5'hf == rd ? _next_reg_rd_12 : _GEN_1036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1069 = 5'h10 == rd ? _next_reg_rd_12 : _GEN_1037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1070 = 5'h11 == rd ? _next_reg_rd_12 : _GEN_1038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1071 = 5'h12 == rd ? _next_reg_rd_12 : _GEN_1039; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1072 = 5'h13 == rd ? _next_reg_rd_12 : _GEN_1040; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1073 = 5'h14 == rd ? _next_reg_rd_12 : _GEN_1041; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1074 = 5'h15 == rd ? _next_reg_rd_12 : _GEN_1042; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1075 = 5'h16 == rd ? _next_reg_rd_12 : _GEN_1043; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1076 = 5'h17 == rd ? _next_reg_rd_12 : _GEN_1044; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1077 = 5'h18 == rd ? _next_reg_rd_12 : _GEN_1045; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1078 = 5'h19 == rd ? _next_reg_rd_12 : _GEN_1046; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1079 = 5'h1a == rd ? _next_reg_rd_12 : _GEN_1047; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1080 = 5'h1b == rd ? _next_reg_rd_12 : _GEN_1048; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1081 = 5'h1c == rd ? _next_reg_rd_12 : _GEN_1049; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1082 = 5'h1d == rd ? _next_reg_rd_12 : _GEN_1050; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1083 = 5'h1e == rd ? _next_reg_rd_12 : _GEN_1051; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1084 = 5'h1f == rd ? _next_reg_rd_12 : _GEN_1052; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:{46,46}]
  wire [63:0] _GEN_1093 = _T_102 ? _GEN_1054 : _GEN_1022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1094 = _T_102 ? _GEN_1055 : _GEN_1023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1095 = _T_102 ? _GEN_1056 : _GEN_1024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1096 = _T_102 ? _GEN_1057 : _GEN_1025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1097 = _T_102 ? _GEN_1058 : _GEN_1026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1098 = _T_102 ? _GEN_1059 : _GEN_1027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1099 = _T_102 ? _GEN_1060 : _GEN_1028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1100 = _T_102 ? _GEN_1061 : _GEN_1029; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1101 = _T_102 ? _GEN_1062 : _GEN_1030; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1102 = _T_102 ? _GEN_1063 : _GEN_1031; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1103 = _T_102 ? _GEN_1064 : _GEN_1032; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1104 = _T_102 ? _GEN_1065 : _GEN_1033; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1105 = _T_102 ? _GEN_1066 : _GEN_1034; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1106 = _T_102 ? _GEN_1067 : _GEN_1035; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1107 = _T_102 ? _GEN_1068 : _GEN_1036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1108 = _T_102 ? _GEN_1069 : _GEN_1037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1109 = _T_102 ? _GEN_1070 : _GEN_1038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1110 = _T_102 ? _GEN_1071 : _GEN_1039; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1111 = _T_102 ? _GEN_1072 : _GEN_1040; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1112 = _T_102 ? _GEN_1073 : _GEN_1041; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1113 = _T_102 ? _GEN_1074 : _GEN_1042; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1114 = _T_102 ? _GEN_1075 : _GEN_1043; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1115 = _T_102 ? _GEN_1076 : _GEN_1044; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1116 = _T_102 ? _GEN_1077 : _GEN_1045; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1117 = _T_102 ? _GEN_1078 : _GEN_1046; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1118 = _T_102 ? _GEN_1079 : _GEN_1047; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1119 = _T_102 ? _GEN_1080 : _GEN_1048; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1120 = _T_102 ? _GEN_1081 : _GEN_1049; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1121 = _T_102 ? _GEN_1082 : _GEN_1050; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1122 = _T_102 ? _GEN_1083 : _GEN_1051; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _GEN_1123 = _T_102 ? _GEN_1084 : _GEN_1052; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 170:22]
  wire [63:0] _next_reg_T_29 = _GEN_101 & _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:61]
  wire [63:0] _GEN_1125 = 5'h1 == rd ? _next_reg_T_29 : _GEN_1093; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1126 = 5'h2 == rd ? _next_reg_T_29 : _GEN_1094; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1127 = 5'h3 == rd ? _next_reg_T_29 : _GEN_1095; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1128 = 5'h4 == rd ? _next_reg_T_29 : _GEN_1096; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1129 = 5'h5 == rd ? _next_reg_T_29 : _GEN_1097; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1130 = 5'h6 == rd ? _next_reg_T_29 : _GEN_1098; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1131 = 5'h7 == rd ? _next_reg_T_29 : _GEN_1099; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1132 = 5'h8 == rd ? _next_reg_T_29 : _GEN_1100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1133 = 5'h9 == rd ? _next_reg_T_29 : _GEN_1101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1134 = 5'ha == rd ? _next_reg_T_29 : _GEN_1102; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1135 = 5'hb == rd ? _next_reg_T_29 : _GEN_1103; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1136 = 5'hc == rd ? _next_reg_T_29 : _GEN_1104; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1137 = 5'hd == rd ? _next_reg_T_29 : _GEN_1105; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1138 = 5'he == rd ? _next_reg_T_29 : _GEN_1106; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1139 = 5'hf == rd ? _next_reg_T_29 : _GEN_1107; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1140 = 5'h10 == rd ? _next_reg_T_29 : _GEN_1108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1141 = 5'h11 == rd ? _next_reg_T_29 : _GEN_1109; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1142 = 5'h12 == rd ? _next_reg_T_29 : _GEN_1110; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1143 = 5'h13 == rd ? _next_reg_T_29 : _GEN_1111; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1144 = 5'h14 == rd ? _next_reg_T_29 : _GEN_1112; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1145 = 5'h15 == rd ? _next_reg_T_29 : _GEN_1113; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1146 = 5'h16 == rd ? _next_reg_T_29 : _GEN_1114; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1147 = 5'h17 == rd ? _next_reg_T_29 : _GEN_1115; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1148 = 5'h18 == rd ? _next_reg_T_29 : _GEN_1116; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1149 = 5'h19 == rd ? _next_reg_T_29 : _GEN_1117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1150 = 5'h1a == rd ? _next_reg_T_29 : _GEN_1118; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1151 = 5'h1b == rd ? _next_reg_T_29 : _GEN_1119; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1152 = 5'h1c == rd ? _next_reg_T_29 : _GEN_1120; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1153 = 5'h1d == rd ? _next_reg_T_29 : _GEN_1121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1154 = 5'h1e == rd ? _next_reg_T_29 : _GEN_1122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1155 = 5'h1f == rd ? _next_reg_T_29 : _GEN_1123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:{45,45}]
  wire [63:0] _GEN_1164 = _T_109 ? _GEN_1125 : _GEN_1093; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1165 = _T_109 ? _GEN_1126 : _GEN_1094; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1166 = _T_109 ? _GEN_1127 : _GEN_1095; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1167 = _T_109 ? _GEN_1128 : _GEN_1096; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1168 = _T_109 ? _GEN_1129 : _GEN_1097; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1169 = _T_109 ? _GEN_1130 : _GEN_1098; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1170 = _T_109 ? _GEN_1131 : _GEN_1099; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1171 = _T_109 ? _GEN_1132 : _GEN_1100; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1172 = _T_109 ? _GEN_1133 : _GEN_1101; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1173 = _T_109 ? _GEN_1134 : _GEN_1102; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1174 = _T_109 ? _GEN_1135 : _GEN_1103; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1175 = _T_109 ? _GEN_1136 : _GEN_1104; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1176 = _T_109 ? _GEN_1137 : _GEN_1105; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1177 = _T_109 ? _GEN_1138 : _GEN_1106; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1178 = _T_109 ? _GEN_1139 : _GEN_1107; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1179 = _T_109 ? _GEN_1140 : _GEN_1108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1180 = _T_109 ? _GEN_1141 : _GEN_1109; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1181 = _T_109 ? _GEN_1142 : _GEN_1110; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1182 = _T_109 ? _GEN_1143 : _GEN_1111; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1183 = _T_109 ? _GEN_1144 : _GEN_1112; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1184 = _T_109 ? _GEN_1145 : _GEN_1113; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1185 = _T_109 ? _GEN_1146 : _GEN_1114; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1186 = _T_109 ? _GEN_1147 : _GEN_1115; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1187 = _T_109 ? _GEN_1148 : _GEN_1116; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1188 = _T_109 ? _GEN_1149 : _GEN_1117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1189 = _T_109 ? _GEN_1150 : _GEN_1118; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1190 = _T_109 ? _GEN_1151 : _GEN_1119; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1191 = _T_109 ? _GEN_1152 : _GEN_1120; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1192 = _T_109 ? _GEN_1153 : _GEN_1121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1193 = _T_109 ? _GEN_1154 : _GEN_1122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _GEN_1194 = _T_109 ? _GEN_1155 : _GEN_1123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 172:21]
  wire [63:0] _next_reg_T_30 = _GEN_101 | _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:61]
  wire [63:0] _GEN_1196 = 5'h1 == rd ? _next_reg_T_30 : _GEN_1164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1197 = 5'h2 == rd ? _next_reg_T_30 : _GEN_1165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1198 = 5'h3 == rd ? _next_reg_T_30 : _GEN_1166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1199 = 5'h4 == rd ? _next_reg_T_30 : _GEN_1167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1200 = 5'h5 == rd ? _next_reg_T_30 : _GEN_1168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1201 = 5'h6 == rd ? _next_reg_T_30 : _GEN_1169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1202 = 5'h7 == rd ? _next_reg_T_30 : _GEN_1170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1203 = 5'h8 == rd ? _next_reg_T_30 : _GEN_1171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1204 = 5'h9 == rd ? _next_reg_T_30 : _GEN_1172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1205 = 5'ha == rd ? _next_reg_T_30 : _GEN_1173; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1206 = 5'hb == rd ? _next_reg_T_30 : _GEN_1174; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1207 = 5'hc == rd ? _next_reg_T_30 : _GEN_1175; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1208 = 5'hd == rd ? _next_reg_T_30 : _GEN_1176; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1209 = 5'he == rd ? _next_reg_T_30 : _GEN_1177; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1210 = 5'hf == rd ? _next_reg_T_30 : _GEN_1178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1211 = 5'h10 == rd ? _next_reg_T_30 : _GEN_1179; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1212 = 5'h11 == rd ? _next_reg_T_30 : _GEN_1180; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1213 = 5'h12 == rd ? _next_reg_T_30 : _GEN_1181; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1214 = 5'h13 == rd ? _next_reg_T_30 : _GEN_1182; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1215 = 5'h14 == rd ? _next_reg_T_30 : _GEN_1183; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1216 = 5'h15 == rd ? _next_reg_T_30 : _GEN_1184; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1217 = 5'h16 == rd ? _next_reg_T_30 : _GEN_1185; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1218 = 5'h17 == rd ? _next_reg_T_30 : _GEN_1186; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1219 = 5'h18 == rd ? _next_reg_T_30 : _GEN_1187; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1220 = 5'h19 == rd ? _next_reg_T_30 : _GEN_1188; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1221 = 5'h1a == rd ? _next_reg_T_30 : _GEN_1189; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1222 = 5'h1b == rd ? _next_reg_T_30 : _GEN_1190; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1223 = 5'h1c == rd ? _next_reg_T_30 : _GEN_1191; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1224 = 5'h1d == rd ? _next_reg_T_30 : _GEN_1192; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1225 = 5'h1e == rd ? _next_reg_T_30 : _GEN_1193; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1226 = 5'h1f == rd ? _next_reg_T_30 : _GEN_1194; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:{45,45}]
  wire [63:0] _GEN_1235 = _T_116 ? _GEN_1196 : _GEN_1164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1236 = _T_116 ? _GEN_1197 : _GEN_1165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1237 = _T_116 ? _GEN_1198 : _GEN_1166; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1238 = _T_116 ? _GEN_1199 : _GEN_1167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1239 = _T_116 ? _GEN_1200 : _GEN_1168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1240 = _T_116 ? _GEN_1201 : _GEN_1169; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1241 = _T_116 ? _GEN_1202 : _GEN_1170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1242 = _T_116 ? _GEN_1203 : _GEN_1171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1243 = _T_116 ? _GEN_1204 : _GEN_1172; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1244 = _T_116 ? _GEN_1205 : _GEN_1173; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1245 = _T_116 ? _GEN_1206 : _GEN_1174; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1246 = _T_116 ? _GEN_1207 : _GEN_1175; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1247 = _T_116 ? _GEN_1208 : _GEN_1176; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1248 = _T_116 ? _GEN_1209 : _GEN_1177; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1249 = _T_116 ? _GEN_1210 : _GEN_1178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1250 = _T_116 ? _GEN_1211 : _GEN_1179; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1251 = _T_116 ? _GEN_1212 : _GEN_1180; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1252 = _T_116 ? _GEN_1213 : _GEN_1181; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1253 = _T_116 ? _GEN_1214 : _GEN_1182; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1254 = _T_116 ? _GEN_1215 : _GEN_1183; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1255 = _T_116 ? _GEN_1216 : _GEN_1184; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1256 = _T_116 ? _GEN_1217 : _GEN_1185; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1257 = _T_116 ? _GEN_1218 : _GEN_1186; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1258 = _T_116 ? _GEN_1219 : _GEN_1187; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1259 = _T_116 ? _GEN_1220 : _GEN_1188; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1260 = _T_116 ? _GEN_1221 : _GEN_1189; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1261 = _T_116 ? _GEN_1222 : _GEN_1190; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1262 = _T_116 ? _GEN_1223 : _GEN_1191; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1263 = _T_116 ? _GEN_1224 : _GEN_1192; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1264 = _T_116 ? _GEN_1225 : _GEN_1193; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _GEN_1265 = _T_116 ? _GEN_1226 : _GEN_1194; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 173:21]
  wire [63:0] _next_reg_T_31 = _GEN_101 ^ _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:61]
  wire [63:0] _GEN_1267 = 5'h1 == rd ? _next_reg_T_31 : _GEN_1235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1268 = 5'h2 == rd ? _next_reg_T_31 : _GEN_1236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1269 = 5'h3 == rd ? _next_reg_T_31 : _GEN_1237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1270 = 5'h4 == rd ? _next_reg_T_31 : _GEN_1238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1271 = 5'h5 == rd ? _next_reg_T_31 : _GEN_1239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1272 = 5'h6 == rd ? _next_reg_T_31 : _GEN_1240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1273 = 5'h7 == rd ? _next_reg_T_31 : _GEN_1241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1274 = 5'h8 == rd ? _next_reg_T_31 : _GEN_1242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1275 = 5'h9 == rd ? _next_reg_T_31 : _GEN_1243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1276 = 5'ha == rd ? _next_reg_T_31 : _GEN_1244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1277 = 5'hb == rd ? _next_reg_T_31 : _GEN_1245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1278 = 5'hc == rd ? _next_reg_T_31 : _GEN_1246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1279 = 5'hd == rd ? _next_reg_T_31 : _GEN_1247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1280 = 5'he == rd ? _next_reg_T_31 : _GEN_1248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1281 = 5'hf == rd ? _next_reg_T_31 : _GEN_1249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1282 = 5'h10 == rd ? _next_reg_T_31 : _GEN_1250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1283 = 5'h11 == rd ? _next_reg_T_31 : _GEN_1251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1284 = 5'h12 == rd ? _next_reg_T_31 : _GEN_1252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1285 = 5'h13 == rd ? _next_reg_T_31 : _GEN_1253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1286 = 5'h14 == rd ? _next_reg_T_31 : _GEN_1254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1287 = 5'h15 == rd ? _next_reg_T_31 : _GEN_1255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1288 = 5'h16 == rd ? _next_reg_T_31 : _GEN_1256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1289 = 5'h17 == rd ? _next_reg_T_31 : _GEN_1257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1290 = 5'h18 == rd ? _next_reg_T_31 : _GEN_1258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1291 = 5'h19 == rd ? _next_reg_T_31 : _GEN_1259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1292 = 5'h1a == rd ? _next_reg_T_31 : _GEN_1260; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1293 = 5'h1b == rd ? _next_reg_T_31 : _GEN_1261; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1294 = 5'h1c == rd ? _next_reg_T_31 : _GEN_1262; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1295 = 5'h1d == rd ? _next_reg_T_31 : _GEN_1263; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1296 = 5'h1e == rd ? _next_reg_T_31 : _GEN_1264; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1297 = 5'h1f == rd ? _next_reg_T_31 : _GEN_1265; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:{45,45}]
  wire [63:0] _GEN_1306 = _T_123 ? _GEN_1267 : _GEN_1235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1307 = _T_123 ? _GEN_1268 : _GEN_1236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1308 = _T_123 ? _GEN_1269 : _GEN_1237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1309 = _T_123 ? _GEN_1270 : _GEN_1238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1310 = _T_123 ? _GEN_1271 : _GEN_1239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1311 = _T_123 ? _GEN_1272 : _GEN_1240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1312 = _T_123 ? _GEN_1273 : _GEN_1241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1313 = _T_123 ? _GEN_1274 : _GEN_1242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1314 = _T_123 ? _GEN_1275 : _GEN_1243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1315 = _T_123 ? _GEN_1276 : _GEN_1244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1316 = _T_123 ? _GEN_1277 : _GEN_1245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1317 = _T_123 ? _GEN_1278 : _GEN_1246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1318 = _T_123 ? _GEN_1279 : _GEN_1247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1319 = _T_123 ? _GEN_1280 : _GEN_1248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1320 = _T_123 ? _GEN_1281 : _GEN_1249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1321 = _T_123 ? _GEN_1282 : _GEN_1250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1322 = _T_123 ? _GEN_1283 : _GEN_1251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1323 = _T_123 ? _GEN_1284 : _GEN_1252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1324 = _T_123 ? _GEN_1285 : _GEN_1253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1325 = _T_123 ? _GEN_1286 : _GEN_1254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1326 = _T_123 ? _GEN_1287 : _GEN_1255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1327 = _T_123 ? _GEN_1288 : _GEN_1256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1328 = _T_123 ? _GEN_1289 : _GEN_1257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1329 = _T_123 ? _GEN_1290 : _GEN_1258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1330 = _T_123 ? _GEN_1291 : _GEN_1259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1331 = _T_123 ? _GEN_1292 : _GEN_1260; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1332 = _T_123 ? _GEN_1293 : _GEN_1261; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1333 = _T_123 ? _GEN_1294 : _GEN_1262; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1334 = _T_123 ? _GEN_1295 : _GEN_1263; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1335 = _T_123 ? _GEN_1296 : _GEN_1264; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [63:0] _GEN_1336 = _T_123 ? _GEN_1297 : _GEN_1265; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 174:21]
  wire [94:0] _GEN_1 = {{31'd0}, _GEN_101}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:61]
  wire [94:0] _next_reg_T_33 = _GEN_1 << _GEN_910[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:61]
  wire [63:0] _GEN_1338 = 5'h1 == rd ? _next_reg_T_33[63:0] : _GEN_1306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1339 = 5'h2 == rd ? _next_reg_T_33[63:0] : _GEN_1307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1340 = 5'h3 == rd ? _next_reg_T_33[63:0] : _GEN_1308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1341 = 5'h4 == rd ? _next_reg_T_33[63:0] : _GEN_1309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1342 = 5'h5 == rd ? _next_reg_T_33[63:0] : _GEN_1310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1343 = 5'h6 == rd ? _next_reg_T_33[63:0] : _GEN_1311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1344 = 5'h7 == rd ? _next_reg_T_33[63:0] : _GEN_1312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1345 = 5'h8 == rd ? _next_reg_T_33[63:0] : _GEN_1313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1346 = 5'h9 == rd ? _next_reg_T_33[63:0] : _GEN_1314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1347 = 5'ha == rd ? _next_reg_T_33[63:0] : _GEN_1315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1348 = 5'hb == rd ? _next_reg_T_33[63:0] : _GEN_1316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1349 = 5'hc == rd ? _next_reg_T_33[63:0] : _GEN_1317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1350 = 5'hd == rd ? _next_reg_T_33[63:0] : _GEN_1318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1351 = 5'he == rd ? _next_reg_T_33[63:0] : _GEN_1319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1352 = 5'hf == rd ? _next_reg_T_33[63:0] : _GEN_1320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1353 = 5'h10 == rd ? _next_reg_T_33[63:0] : _GEN_1321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1354 = 5'h11 == rd ? _next_reg_T_33[63:0] : _GEN_1322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1355 = 5'h12 == rd ? _next_reg_T_33[63:0] : _GEN_1323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1356 = 5'h13 == rd ? _next_reg_T_33[63:0] : _GEN_1324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1357 = 5'h14 == rd ? _next_reg_T_33[63:0] : _GEN_1325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1358 = 5'h15 == rd ? _next_reg_T_33[63:0] : _GEN_1326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1359 = 5'h16 == rd ? _next_reg_T_33[63:0] : _GEN_1327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1360 = 5'h17 == rd ? _next_reg_T_33[63:0] : _GEN_1328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1361 = 5'h18 == rd ? _next_reg_T_33[63:0] : _GEN_1329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1362 = 5'h19 == rd ? _next_reg_T_33[63:0] : _GEN_1330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1363 = 5'h1a == rd ? _next_reg_T_33[63:0] : _GEN_1331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1364 = 5'h1b == rd ? _next_reg_T_33[63:0] : _GEN_1332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1365 = 5'h1c == rd ? _next_reg_T_33[63:0] : _GEN_1333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1366 = 5'h1d == rd ? _next_reg_T_33[63:0] : _GEN_1334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1367 = 5'h1e == rd ? _next_reg_T_33[63:0] : _GEN_1335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1368 = 5'h1f == rd ? _next_reg_T_33[63:0] : _GEN_1336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:{45,45}]
  wire [63:0] _GEN_1377 = _T_762 ? _GEN_1338 : _GEN_1306; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1378 = _T_762 ? _GEN_1339 : _GEN_1307; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1379 = _T_762 ? _GEN_1340 : _GEN_1308; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1380 = _T_762 ? _GEN_1341 : _GEN_1309; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1381 = _T_762 ? _GEN_1342 : _GEN_1310; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1382 = _T_762 ? _GEN_1343 : _GEN_1311; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1383 = _T_762 ? _GEN_1344 : _GEN_1312; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1384 = _T_762 ? _GEN_1345 : _GEN_1313; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1385 = _T_762 ? _GEN_1346 : _GEN_1314; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1386 = _T_762 ? _GEN_1347 : _GEN_1315; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1387 = _T_762 ? _GEN_1348 : _GEN_1316; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1388 = _T_762 ? _GEN_1349 : _GEN_1317; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1389 = _T_762 ? _GEN_1350 : _GEN_1318; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1390 = _T_762 ? _GEN_1351 : _GEN_1319; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1391 = _T_762 ? _GEN_1352 : _GEN_1320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1392 = _T_762 ? _GEN_1353 : _GEN_1321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1393 = _T_762 ? _GEN_1354 : _GEN_1322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1394 = _T_762 ? _GEN_1355 : _GEN_1323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1395 = _T_762 ? _GEN_1356 : _GEN_1324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1396 = _T_762 ? _GEN_1357 : _GEN_1325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1397 = _T_762 ? _GEN_1358 : _GEN_1326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1398 = _T_762 ? _GEN_1359 : _GEN_1327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1399 = _T_762 ? _GEN_1360 : _GEN_1328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1400 = _T_762 ? _GEN_1361 : _GEN_1329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1401 = _T_762 ? _GEN_1362 : _GEN_1330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1402 = _T_762 ? _GEN_1363 : _GEN_1331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1403 = _T_762 ? _GEN_1364 : _GEN_1332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1404 = _T_762 ? _GEN_1365 : _GEN_1333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1405 = _T_762 ? _GEN_1366 : _GEN_1334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1406 = _T_762 ? _GEN_1367 : _GEN_1335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _GEN_1407 = _T_762 ? _GEN_1368 : _GEN_1336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 176:21]
  wire [63:0] _next_reg_T_35 = _GEN_101 >> _GEN_910[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:61]
  wire [63:0] _GEN_1409 = 5'h1 == rd ? _next_reg_T_35 : _GEN_1377; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1410 = 5'h2 == rd ? _next_reg_T_35 : _GEN_1378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1411 = 5'h3 == rd ? _next_reg_T_35 : _GEN_1379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1412 = 5'h4 == rd ? _next_reg_T_35 : _GEN_1380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1413 = 5'h5 == rd ? _next_reg_T_35 : _GEN_1381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1414 = 5'h6 == rd ? _next_reg_T_35 : _GEN_1382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1415 = 5'h7 == rd ? _next_reg_T_35 : _GEN_1383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1416 = 5'h8 == rd ? _next_reg_T_35 : _GEN_1384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1417 = 5'h9 == rd ? _next_reg_T_35 : _GEN_1385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1418 = 5'ha == rd ? _next_reg_T_35 : _GEN_1386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1419 = 5'hb == rd ? _next_reg_T_35 : _GEN_1387; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1420 = 5'hc == rd ? _next_reg_T_35 : _GEN_1388; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1421 = 5'hd == rd ? _next_reg_T_35 : _GEN_1389; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1422 = 5'he == rd ? _next_reg_T_35 : _GEN_1390; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1423 = 5'hf == rd ? _next_reg_T_35 : _GEN_1391; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1424 = 5'h10 == rd ? _next_reg_T_35 : _GEN_1392; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1425 = 5'h11 == rd ? _next_reg_T_35 : _GEN_1393; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1426 = 5'h12 == rd ? _next_reg_T_35 : _GEN_1394; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1427 = 5'h13 == rd ? _next_reg_T_35 : _GEN_1395; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1428 = 5'h14 == rd ? _next_reg_T_35 : _GEN_1396; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1429 = 5'h15 == rd ? _next_reg_T_35 : _GEN_1397; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1430 = 5'h16 == rd ? _next_reg_T_35 : _GEN_1398; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1431 = 5'h17 == rd ? _next_reg_T_35 : _GEN_1399; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1432 = 5'h18 == rd ? _next_reg_T_35 : _GEN_1400; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1433 = 5'h19 == rd ? _next_reg_T_35 : _GEN_1401; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1434 = 5'h1a == rd ? _next_reg_T_35 : _GEN_1402; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1435 = 5'h1b == rd ? _next_reg_T_35 : _GEN_1403; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1436 = 5'h1c == rd ? _next_reg_T_35 : _GEN_1404; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1437 = 5'h1d == rd ? _next_reg_T_35 : _GEN_1405; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1438 = 5'h1e == rd ? _next_reg_T_35 : _GEN_1406; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1439 = 5'h1f == rd ? _next_reg_T_35 : _GEN_1407; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:{45,45}]
  wire [63:0] _GEN_1448 = _T_769 ? _GEN_1409 : _GEN_1377; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1449 = _T_769 ? _GEN_1410 : _GEN_1378; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1450 = _T_769 ? _GEN_1411 : _GEN_1379; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1451 = _T_769 ? _GEN_1412 : _GEN_1380; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1452 = _T_769 ? _GEN_1413 : _GEN_1381; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1453 = _T_769 ? _GEN_1414 : _GEN_1382; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1454 = _T_769 ? _GEN_1415 : _GEN_1383; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1455 = _T_769 ? _GEN_1416 : _GEN_1384; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1456 = _T_769 ? _GEN_1417 : _GEN_1385; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1457 = _T_769 ? _GEN_1418 : _GEN_1386; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1458 = _T_769 ? _GEN_1419 : _GEN_1387; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1459 = _T_769 ? _GEN_1420 : _GEN_1388; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1460 = _T_769 ? _GEN_1421 : _GEN_1389; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1461 = _T_769 ? _GEN_1422 : _GEN_1390; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1462 = _T_769 ? _GEN_1423 : _GEN_1391; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1463 = _T_769 ? _GEN_1424 : _GEN_1392; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1464 = _T_769 ? _GEN_1425 : _GEN_1393; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1465 = _T_769 ? _GEN_1426 : _GEN_1394; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1466 = _T_769 ? _GEN_1427 : _GEN_1395; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1467 = _T_769 ? _GEN_1428 : _GEN_1396; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1468 = _T_769 ? _GEN_1429 : _GEN_1397; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1469 = _T_769 ? _GEN_1430 : _GEN_1398; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1470 = _T_769 ? _GEN_1431 : _GEN_1399; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1471 = _T_769 ? _GEN_1432 : _GEN_1400; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1472 = _T_769 ? _GEN_1433 : _GEN_1401; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1473 = _T_769 ? _GEN_1434 : _GEN_1402; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1474 = _T_769 ? _GEN_1435 : _GEN_1403; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1475 = _T_769 ? _GEN_1436 : _GEN_1404; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1476 = _T_769 ? _GEN_1437 : _GEN_1405; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1477 = _T_769 ? _GEN_1438 : _GEN_1406; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _GEN_1478 = _T_769 ? _GEN_1439 : _GEN_1407; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 177:21]
  wire [63:0] _next_reg_T_37 = _GEN_101 - _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:61]
  wire [63:0] _GEN_1480 = 5'h1 == rd ? _next_reg_T_37 : _GEN_1448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1481 = 5'h2 == rd ? _next_reg_T_37 : _GEN_1449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1482 = 5'h3 == rd ? _next_reg_T_37 : _GEN_1450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1483 = 5'h4 == rd ? _next_reg_T_37 : _GEN_1451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1484 = 5'h5 == rd ? _next_reg_T_37 : _GEN_1452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1485 = 5'h6 == rd ? _next_reg_T_37 : _GEN_1453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1486 = 5'h7 == rd ? _next_reg_T_37 : _GEN_1454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1487 = 5'h8 == rd ? _next_reg_T_37 : _GEN_1455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1488 = 5'h9 == rd ? _next_reg_T_37 : _GEN_1456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1489 = 5'ha == rd ? _next_reg_T_37 : _GEN_1457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1490 = 5'hb == rd ? _next_reg_T_37 : _GEN_1458; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1491 = 5'hc == rd ? _next_reg_T_37 : _GEN_1459; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1492 = 5'hd == rd ? _next_reg_T_37 : _GEN_1460; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1493 = 5'he == rd ? _next_reg_T_37 : _GEN_1461; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1494 = 5'hf == rd ? _next_reg_T_37 : _GEN_1462; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1495 = 5'h10 == rd ? _next_reg_T_37 : _GEN_1463; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1496 = 5'h11 == rd ? _next_reg_T_37 : _GEN_1464; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1497 = 5'h12 == rd ? _next_reg_T_37 : _GEN_1465; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1498 = 5'h13 == rd ? _next_reg_T_37 : _GEN_1466; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1499 = 5'h14 == rd ? _next_reg_T_37 : _GEN_1467; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1500 = 5'h15 == rd ? _next_reg_T_37 : _GEN_1468; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1501 = 5'h16 == rd ? _next_reg_T_37 : _GEN_1469; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1502 = 5'h17 == rd ? _next_reg_T_37 : _GEN_1470; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1503 = 5'h18 == rd ? _next_reg_T_37 : _GEN_1471; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1504 = 5'h19 == rd ? _next_reg_T_37 : _GEN_1472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1505 = 5'h1a == rd ? _next_reg_T_37 : _GEN_1473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1506 = 5'h1b == rd ? _next_reg_T_37 : _GEN_1474; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1507 = 5'h1c == rd ? _next_reg_T_37 : _GEN_1475; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1508 = 5'h1d == rd ? _next_reg_T_37 : _GEN_1476; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1509 = 5'h1e == rd ? _next_reg_T_37 : _GEN_1477; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1510 = 5'h1f == rd ? _next_reg_T_37 : _GEN_1478; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:{45,45}]
  wire [63:0] _GEN_1519 = _T_144 ? _GEN_1480 : _GEN_1448; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1520 = _T_144 ? _GEN_1481 : _GEN_1449; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1521 = _T_144 ? _GEN_1482 : _GEN_1450; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1522 = _T_144 ? _GEN_1483 : _GEN_1451; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1523 = _T_144 ? _GEN_1484 : _GEN_1452; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1524 = _T_144 ? _GEN_1485 : _GEN_1453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1525 = _T_144 ? _GEN_1486 : _GEN_1454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1526 = _T_144 ? _GEN_1487 : _GEN_1455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1527 = _T_144 ? _GEN_1488 : _GEN_1456; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1528 = _T_144 ? _GEN_1489 : _GEN_1457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1529 = _T_144 ? _GEN_1490 : _GEN_1458; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1530 = _T_144 ? _GEN_1491 : _GEN_1459; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1531 = _T_144 ? _GEN_1492 : _GEN_1460; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1532 = _T_144 ? _GEN_1493 : _GEN_1461; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1533 = _T_144 ? _GEN_1494 : _GEN_1462; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1534 = _T_144 ? _GEN_1495 : _GEN_1463; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1535 = _T_144 ? _GEN_1496 : _GEN_1464; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1536 = _T_144 ? _GEN_1497 : _GEN_1465; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1537 = _T_144 ? _GEN_1498 : _GEN_1466; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1538 = _T_144 ? _GEN_1499 : _GEN_1467; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1539 = _T_144 ? _GEN_1500 : _GEN_1468; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1540 = _T_144 ? _GEN_1501 : _GEN_1469; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1541 = _T_144 ? _GEN_1502 : _GEN_1470; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1542 = _T_144 ? _GEN_1503 : _GEN_1471; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1543 = _T_144 ? _GEN_1504 : _GEN_1472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1544 = _T_144 ? _GEN_1505 : _GEN_1473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1545 = _T_144 ? _GEN_1506 : _GEN_1474; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1546 = _T_144 ? _GEN_1507 : _GEN_1475; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1547 = _T_144 ? _GEN_1508 : _GEN_1476; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1548 = _T_144 ? _GEN_1509 : _GEN_1477; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _GEN_1549 = _T_144 ? _GEN_1510 : _GEN_1478; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 179:21]
  wire [63:0] _next_reg_T_41 = $signed(_T_325) >>> _GEN_910[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:92]
  wire [63:0] _GEN_1551 = 5'h1 == rd ? _next_reg_T_41 : _GEN_1519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1552 = 5'h2 == rd ? _next_reg_T_41 : _GEN_1520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1553 = 5'h3 == rd ? _next_reg_T_41 : _GEN_1521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1554 = 5'h4 == rd ? _next_reg_T_41 : _GEN_1522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1555 = 5'h5 == rd ? _next_reg_T_41 : _GEN_1523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1556 = 5'h6 == rd ? _next_reg_T_41 : _GEN_1524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1557 = 5'h7 == rd ? _next_reg_T_41 : _GEN_1525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1558 = 5'h8 == rd ? _next_reg_T_41 : _GEN_1526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1559 = 5'h9 == rd ? _next_reg_T_41 : _GEN_1527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1560 = 5'ha == rd ? _next_reg_T_41 : _GEN_1528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1561 = 5'hb == rd ? _next_reg_T_41 : _GEN_1529; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1562 = 5'hc == rd ? _next_reg_T_41 : _GEN_1530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1563 = 5'hd == rd ? _next_reg_T_41 : _GEN_1531; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1564 = 5'he == rd ? _next_reg_T_41 : _GEN_1532; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1565 = 5'hf == rd ? _next_reg_T_41 : _GEN_1533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1566 = 5'h10 == rd ? _next_reg_T_41 : _GEN_1534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1567 = 5'h11 == rd ? _next_reg_T_41 : _GEN_1535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1568 = 5'h12 == rd ? _next_reg_T_41 : _GEN_1536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1569 = 5'h13 == rd ? _next_reg_T_41 : _GEN_1537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1570 = 5'h14 == rd ? _next_reg_T_41 : _GEN_1538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1571 = 5'h15 == rd ? _next_reg_T_41 : _GEN_1539; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1572 = 5'h16 == rd ? _next_reg_T_41 : _GEN_1540; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1573 = 5'h17 == rd ? _next_reg_T_41 : _GEN_1541; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1574 = 5'h18 == rd ? _next_reg_T_41 : _GEN_1542; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1575 = 5'h19 == rd ? _next_reg_T_41 : _GEN_1543; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1576 = 5'h1a == rd ? _next_reg_T_41 : _GEN_1544; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1577 = 5'h1b == rd ? _next_reg_T_41 : _GEN_1545; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1578 = 5'h1c == rd ? _next_reg_T_41 : _GEN_1546; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1579 = 5'h1d == rd ? _next_reg_T_41 : _GEN_1547; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1580 = 5'h1e == rd ? _next_reg_T_41 : _GEN_1548; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1581 = 5'h1f == rd ? _next_reg_T_41 : _GEN_1549; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:{45,45}]
  wire [63:0] _GEN_1590 = _T_776 ? _GEN_1551 : _GEN_1519; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1591 = _T_776 ? _GEN_1552 : _GEN_1520; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1592 = _T_776 ? _GEN_1553 : _GEN_1521; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1593 = _T_776 ? _GEN_1554 : _GEN_1522; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1594 = _T_776 ? _GEN_1555 : _GEN_1523; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1595 = _T_776 ? _GEN_1556 : _GEN_1524; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1596 = _T_776 ? _GEN_1557 : _GEN_1525; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1597 = _T_776 ? _GEN_1558 : _GEN_1526; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1598 = _T_776 ? _GEN_1559 : _GEN_1527; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1599 = _T_776 ? _GEN_1560 : _GEN_1528; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1600 = _T_776 ? _GEN_1561 : _GEN_1529; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1601 = _T_776 ? _GEN_1562 : _GEN_1530; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1602 = _T_776 ? _GEN_1563 : _GEN_1531; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1603 = _T_776 ? _GEN_1564 : _GEN_1532; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1604 = _T_776 ? _GEN_1565 : _GEN_1533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1605 = _T_776 ? _GEN_1566 : _GEN_1534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1606 = _T_776 ? _GEN_1567 : _GEN_1535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1607 = _T_776 ? _GEN_1568 : _GEN_1536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1608 = _T_776 ? _GEN_1569 : _GEN_1537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1609 = _T_776 ? _GEN_1570 : _GEN_1538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1610 = _T_776 ? _GEN_1571 : _GEN_1539; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1611 = _T_776 ? _GEN_1572 : _GEN_1540; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1612 = _T_776 ? _GEN_1573 : _GEN_1541; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1613 = _T_776 ? _GEN_1574 : _GEN_1542; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1614 = _T_776 ? _GEN_1575 : _GEN_1543; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1615 = _T_776 ? _GEN_1576 : _GEN_1544; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1616 = _T_776 ? _GEN_1577 : _GEN_1545; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1617 = _T_776 ? _GEN_1578 : _GEN_1546; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1618 = _T_776 ? _GEN_1579 : _GEN_1547; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1619 = _T_776 ? _GEN_1580 : _GEN_1548; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _GEN_1620 = _T_776 ? _GEN_1581 : _GEN_1549; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 180:21]
  wire [63:0] _next_reg_T_43 = io_now_pc + 64'h4; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:37]
  wire [63:0] _GEN_1622 = 5'h1 == rd ? _next_reg_T_43 : _GEN_1590; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1623 = 5'h2 == rd ? _next_reg_T_43 : _GEN_1591; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1624 = 5'h3 == rd ? _next_reg_T_43 : _GEN_1592; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1625 = 5'h4 == rd ? _next_reg_T_43 : _GEN_1593; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1626 = 5'h5 == rd ? _next_reg_T_43 : _GEN_1594; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1627 = 5'h6 == rd ? _next_reg_T_43 : _GEN_1595; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1628 = 5'h7 == rd ? _next_reg_T_43 : _GEN_1596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1629 = 5'h8 == rd ? _next_reg_T_43 : _GEN_1597; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1630 = 5'h9 == rd ? _next_reg_T_43 : _GEN_1598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1631 = 5'ha == rd ? _next_reg_T_43 : _GEN_1599; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1632 = 5'hb == rd ? _next_reg_T_43 : _GEN_1600; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1633 = 5'hc == rd ? _next_reg_T_43 : _GEN_1601; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1634 = 5'hd == rd ? _next_reg_T_43 : _GEN_1602; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1635 = 5'he == rd ? _next_reg_T_43 : _GEN_1603; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1636 = 5'hf == rd ? _next_reg_T_43 : _GEN_1604; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1637 = 5'h10 == rd ? _next_reg_T_43 : _GEN_1605; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1638 = 5'h11 == rd ? _next_reg_T_43 : _GEN_1606; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1639 = 5'h12 == rd ? _next_reg_T_43 : _GEN_1607; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1640 = 5'h13 == rd ? _next_reg_T_43 : _GEN_1608; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1641 = 5'h14 == rd ? _next_reg_T_43 : _GEN_1609; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1642 = 5'h15 == rd ? _next_reg_T_43 : _GEN_1610; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1643 = 5'h16 == rd ? _next_reg_T_43 : _GEN_1611; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1644 = 5'h17 == rd ? _next_reg_T_43 : _GEN_1612; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1645 = 5'h18 == rd ? _next_reg_T_43 : _GEN_1613; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1646 = 5'h19 == rd ? _next_reg_T_43 : _GEN_1614; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1647 = 5'h1a == rd ? _next_reg_T_43 : _GEN_1615; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1648 = 5'h1b == rd ? _next_reg_T_43 : _GEN_1616; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1649 = 5'h1c == rd ? _next_reg_T_43 : _GEN_1617; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1650 = 5'h1d == rd ? _next_reg_T_43 : _GEN_1618; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1651 = 5'h1e == rd ? _next_reg_T_43 : _GEN_1619; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1652 = 5'h1f == rd ? _next_reg_T_43 : _GEN_1620; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 192:{27,27}]
  wire [63:0] _GEN_1654 = _T_371 ? _T_359 : io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55 191:27]
  wire [63:0] _GEN_1656 = _T_371 ? _GEN_1622 : _GEN_1590; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1657 = _T_371 ? _GEN_1623 : _GEN_1591; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1658 = _T_371 ? _GEN_1624 : _GEN_1592; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1659 = _T_371 ? _GEN_1625 : _GEN_1593; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1660 = _T_371 ? _GEN_1626 : _GEN_1594; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1661 = _T_371 ? _GEN_1627 : _GEN_1595; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1662 = _T_371 ? _GEN_1628 : _GEN_1596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1663 = _T_371 ? _GEN_1629 : _GEN_1597; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1664 = _T_371 ? _GEN_1630 : _GEN_1598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1665 = _T_371 ? _GEN_1631 : _GEN_1599; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1666 = _T_371 ? _GEN_1632 : _GEN_1600; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1667 = _T_371 ? _GEN_1633 : _GEN_1601; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1668 = _T_371 ? _GEN_1634 : _GEN_1602; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1669 = _T_371 ? _GEN_1635 : _GEN_1603; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1670 = _T_371 ? _GEN_1636 : _GEN_1604; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1671 = _T_371 ? _GEN_1637 : _GEN_1605; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1672 = _T_371 ? _GEN_1638 : _GEN_1606; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1673 = _T_371 ? _GEN_1639 : _GEN_1607; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1674 = _T_371 ? _GEN_1640 : _GEN_1608; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1675 = _T_371 ? _GEN_1641 : _GEN_1609; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1676 = _T_371 ? _GEN_1642 : _GEN_1610; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1677 = _T_371 ? _GEN_1643 : _GEN_1611; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1678 = _T_371 ? _GEN_1644 : _GEN_1612; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1679 = _T_371 ? _GEN_1645 : _GEN_1613; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1680 = _T_371 ? _GEN_1646 : _GEN_1614; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1681 = _T_371 ? _GEN_1647 : _GEN_1615; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1682 = _T_371 ? _GEN_1648 : _GEN_1616; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1683 = _T_371 ? _GEN_1649 : _GEN_1617; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1684 = _T_371 ? _GEN_1650 : _GEN_1618; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1685 = _T_371 ? _GEN_1651 : _GEN_1619; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1686 = _T_371 ? _GEN_1652 : _GEN_1620; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55]
  wire [63:0] _GEN_1687 = _T_371 ? io_now_csr_mtval : _T_359; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55 194:24]
  wire  _GEN_1689 = _T_371 ? vmEnable : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 189:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1698 = _T_158 & _T_371; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 113:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1699 = _T_158 ? _GEN_1654 : io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1701 = _T_158 ? _GEN_1656 : _GEN_1590; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1702 = _T_158 ? _GEN_1657 : _GEN_1591; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1703 = _T_158 ? _GEN_1658 : _GEN_1592; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1704 = _T_158 ? _GEN_1659 : _GEN_1593; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1705 = _T_158 ? _GEN_1660 : _GEN_1594; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1706 = _T_158 ? _GEN_1661 : _GEN_1595; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1707 = _T_158 ? _GEN_1662 : _GEN_1596; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1708 = _T_158 ? _GEN_1663 : _GEN_1597; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1709 = _T_158 ? _GEN_1664 : _GEN_1598; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1710 = _T_158 ? _GEN_1665 : _GEN_1599; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1711 = _T_158 ? _GEN_1666 : _GEN_1600; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1712 = _T_158 ? _GEN_1667 : _GEN_1601; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1713 = _T_158 ? _GEN_1668 : _GEN_1602; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1714 = _T_158 ? _GEN_1669 : _GEN_1603; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1715 = _T_158 ? _GEN_1670 : _GEN_1604; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1716 = _T_158 ? _GEN_1671 : _GEN_1605; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1717 = _T_158 ? _GEN_1672 : _GEN_1606; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1718 = _T_158 ? _GEN_1673 : _GEN_1607; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1719 = _T_158 ? _GEN_1674 : _GEN_1608; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1720 = _T_158 ? _GEN_1675 : _GEN_1609; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1721 = _T_158 ? _GEN_1676 : _GEN_1610; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1722 = _T_158 ? _GEN_1677 : _GEN_1611; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1723 = _T_158 ? _GEN_1678 : _GEN_1612; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1724 = _T_158 ? _GEN_1679 : _GEN_1613; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1725 = _T_158 ? _GEN_1680 : _GEN_1614; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1726 = _T_158 ? _GEN_1681 : _GEN_1615; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1727 = _T_158 ? _GEN_1682 : _GEN_1616; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1728 = _T_158 ? _GEN_1683 : _GEN_1617; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1729 = _T_158 ? _GEN_1684 : _GEN_1618; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1730 = _T_158 ? _GEN_1685 : _GEN_1619; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1731 = _T_158 ? _GEN_1686 : _GEN_1620; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1732 = _T_158 ? _GEN_1687 : io_now_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire  _GEN_1734 = _T_158 ? _GEN_1689 : vmEnable; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 187:21]
  wire [63:0] _GEN_1736 = 5'h1 == rd ? _next_reg_T_43 : _GEN_1701; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1737 = 5'h2 == rd ? _next_reg_T_43 : _GEN_1702; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1738 = 5'h3 == rd ? _next_reg_T_43 : _GEN_1703; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1739 = 5'h4 == rd ? _next_reg_T_43 : _GEN_1704; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1740 = 5'h5 == rd ? _next_reg_T_43 : _GEN_1705; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1741 = 5'h6 == rd ? _next_reg_T_43 : _GEN_1706; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1742 = 5'h7 == rd ? _next_reg_T_43 : _GEN_1707; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1743 = 5'h8 == rd ? _next_reg_T_43 : _GEN_1708; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1744 = 5'h9 == rd ? _next_reg_T_43 : _GEN_1709; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1745 = 5'ha == rd ? _next_reg_T_43 : _GEN_1710; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1746 = 5'hb == rd ? _next_reg_T_43 : _GEN_1711; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1747 = 5'hc == rd ? _next_reg_T_43 : _GEN_1712; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1748 = 5'hd == rd ? _next_reg_T_43 : _GEN_1713; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1749 = 5'he == rd ? _next_reg_T_43 : _GEN_1714; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1750 = 5'hf == rd ? _next_reg_T_43 : _GEN_1715; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1751 = 5'h10 == rd ? _next_reg_T_43 : _GEN_1716; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1752 = 5'h11 == rd ? _next_reg_T_43 : _GEN_1717; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1753 = 5'h12 == rd ? _next_reg_T_43 : _GEN_1718; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1754 = 5'h13 == rd ? _next_reg_T_43 : _GEN_1719; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1755 = 5'h14 == rd ? _next_reg_T_43 : _GEN_1720; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1756 = 5'h15 == rd ? _next_reg_T_43 : _GEN_1721; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1757 = 5'h16 == rd ? _next_reg_T_43 : _GEN_1722; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1758 = 5'h17 == rd ? _next_reg_T_43 : _GEN_1723; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1759 = 5'h18 == rd ? _next_reg_T_43 : _GEN_1724; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1760 = 5'h19 == rd ? _next_reg_T_43 : _GEN_1725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1761 = 5'h1a == rd ? _next_reg_T_43 : _GEN_1726; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1762 = 5'h1b == rd ? _next_reg_T_43 : _GEN_1727; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1763 = 5'h1c == rd ? _next_reg_T_43 : _GEN_1728; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1764 = 5'h1d == rd ? _next_reg_T_43 : _GEN_1729; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1765 = 5'h1e == rd ? _next_reg_T_43 : _GEN_1730; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire [63:0] _GEN_1766 = 5'h1f == rd ? _next_reg_T_43 : _GEN_1731; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 204:{27,27}]
  wire  _GEN_1767 = _T_205 | _GEN_1698; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 202:27]
  wire [63:0] _GEN_1768 = _T_205 ? _T_193 : _GEN_1699; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 203:27]
  wire [63:0] _GEN_1770 = _T_205 ? _GEN_1736 : _GEN_1701; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1771 = _T_205 ? _GEN_1737 : _GEN_1702; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1772 = _T_205 ? _GEN_1738 : _GEN_1703; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1773 = _T_205 ? _GEN_1739 : _GEN_1704; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1774 = _T_205 ? _GEN_1740 : _GEN_1705; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1775 = _T_205 ? _GEN_1741 : _GEN_1706; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1776 = _T_205 ? _GEN_1742 : _GEN_1707; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1777 = _T_205 ? _GEN_1743 : _GEN_1708; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1778 = _T_205 ? _GEN_1744 : _GEN_1709; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1779 = _T_205 ? _GEN_1745 : _GEN_1710; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1780 = _T_205 ? _GEN_1746 : _GEN_1711; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1781 = _T_205 ? _GEN_1747 : _GEN_1712; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1782 = _T_205 ? _GEN_1748 : _GEN_1713; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1783 = _T_205 ? _GEN_1749 : _GEN_1714; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1784 = _T_205 ? _GEN_1750 : _GEN_1715; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1785 = _T_205 ? _GEN_1751 : _GEN_1716; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1786 = _T_205 ? _GEN_1752 : _GEN_1717; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1787 = _T_205 ? _GEN_1753 : _GEN_1718; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1788 = _T_205 ? _GEN_1754 : _GEN_1719; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1789 = _T_205 ? _GEN_1755 : _GEN_1720; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1790 = _T_205 ? _GEN_1756 : _GEN_1721; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1791 = _T_205 ? _GEN_1757 : _GEN_1722; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1792 = _T_205 ? _GEN_1758 : _GEN_1723; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1793 = _T_205 ? _GEN_1759 : _GEN_1724; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1794 = _T_205 ? _GEN_1760 : _GEN_1725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1795 = _T_205 ? _GEN_1761 : _GEN_1726; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1796 = _T_205 ? _GEN_1762 : _GEN_1727; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1797 = _T_205 ? _GEN_1763 : _GEN_1728; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1798 = _T_205 ? _GEN_1764 : _GEN_1729; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1799 = _T_205 ? _GEN_1765 : _GEN_1730; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1800 = _T_205 ? _GEN_1766 : _GEN_1731; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91]
  wire [63:0] _GEN_1801 = _T_205 ? _GEN_1732 : _T_193; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 206:24]
  wire  _GEN_1803 = _T_205 ? _GEN_1734 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 201:91 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1811 = _T_182 ? _GEN_1767 : _GEN_1698; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1812 = _T_182 ? _GEN_1768 : _GEN_1699; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1814 = _T_182 ? _GEN_1770 : _GEN_1701; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1815 = _T_182 ? _GEN_1771 : _GEN_1702; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1816 = _T_182 ? _GEN_1772 : _GEN_1703; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1817 = _T_182 ? _GEN_1773 : _GEN_1704; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1818 = _T_182 ? _GEN_1774 : _GEN_1705; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1819 = _T_182 ? _GEN_1775 : _GEN_1706; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1820 = _T_182 ? _GEN_1776 : _GEN_1707; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1821 = _T_182 ? _GEN_1777 : _GEN_1708; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1822 = _T_182 ? _GEN_1778 : _GEN_1709; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1823 = _T_182 ? _GEN_1779 : _GEN_1710; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1824 = _T_182 ? _GEN_1780 : _GEN_1711; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1825 = _T_182 ? _GEN_1781 : _GEN_1712; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1826 = _T_182 ? _GEN_1782 : _GEN_1713; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1827 = _T_182 ? _GEN_1783 : _GEN_1714; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1828 = _T_182 ? _GEN_1784 : _GEN_1715; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1829 = _T_182 ? _GEN_1785 : _GEN_1716; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1830 = _T_182 ? _GEN_1786 : _GEN_1717; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1831 = _T_182 ? _GEN_1787 : _GEN_1718; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1832 = _T_182 ? _GEN_1788 : _GEN_1719; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1833 = _T_182 ? _GEN_1789 : _GEN_1720; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1834 = _T_182 ? _GEN_1790 : _GEN_1721; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1835 = _T_182 ? _GEN_1791 : _GEN_1722; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1836 = _T_182 ? _GEN_1792 : _GEN_1723; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1837 = _T_182 ? _GEN_1793 : _GEN_1724; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1838 = _T_182 ? _GEN_1794 : _GEN_1725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1839 = _T_182 ? _GEN_1795 : _GEN_1726; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1840 = _T_182 ? _GEN_1796 : _GEN_1727; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1841 = _T_182 ? _GEN_1797 : _GEN_1728; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1842 = _T_182 ? _GEN_1798 : _GEN_1729; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1843 = _T_182 ? _GEN_1799 : _GEN_1730; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1844 = _T_182 ? _GEN_1800 : _GEN_1731; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire [63:0] _GEN_1845 = _T_182 ? _GEN_1801 : _GEN_1732; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire  _GEN_1847 = _T_182 ? _GEN_1803 : _GEN_1734; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 199:22]
  wire  _GEN_1848 = _T_371 | _GEN_1811; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 216:29]
  wire [63:0] _GEN_1849 = _T_371 ? _T_359 : _GEN_1812; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 217:29]
  wire [63:0] _GEN_1850 = _T_371 ? _GEN_1845 : _T_359; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 219:26]
  wire  _GEN_1852 = _T_371 ? _GEN_1847 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 215:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1853 = _GEN_101 == _GEN_910 ? _GEN_1848 : _GEN_1811; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire [63:0] _GEN_1854 = _GEN_101 == _GEN_910 ? _GEN_1849 : _GEN_1812; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire [63:0] _GEN_1855 = _GEN_101 == _GEN_910 ? _GEN_1850 : _GEN_1845; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire  _GEN_1857 = _GEN_101 == _GEN_910 ? _GEN_1852 : _GEN_1847; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 214:43]
  wire  _GEN_1868 = _T_207 ? _GEN_1853 : _GEN_1811; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire [63:0] _GEN_1869 = _T_207 ? _GEN_1854 : _GEN_1812; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire [63:0] _GEN_1870 = _T_207 ? _GEN_1855 : _GEN_1845; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire  _GEN_1872 = _T_207 ? _GEN_1857 : _GEN_1847; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 212:21]
  wire  _GEN_1873 = _T_371 | _GEN_1868; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 228:29]
  wire [63:0] _GEN_1874 = _T_371 ? _T_359 : _GEN_1869; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 229:29]
  wire [63:0] _GEN_1875 = _T_371 ? _GEN_1870 : _T_359; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 231:26]
  wire  _GEN_1877 = _T_371 ? _GEN_1872 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 227:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1878 = _GEN_101 != _GEN_910 ? _GEN_1873 : _GEN_1868; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire [63:0] _GEN_1879 = _GEN_101 != _GEN_910 ? _GEN_1874 : _GEN_1869; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire [63:0] _GEN_1880 = _GEN_101 != _GEN_910 ? _GEN_1875 : _GEN_1870; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire  _GEN_1882 = _GEN_101 != _GEN_910 ? _GEN_1877 : _GEN_1872; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 226:43]
  wire  _GEN_1893 = _T_234 ? _GEN_1878 : _GEN_1868; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire [63:0] _GEN_1894 = _T_234 ? _GEN_1879 : _GEN_1869; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire [63:0] _GEN_1895 = _T_234 ? _GEN_1880 : _GEN_1870; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire  _GEN_1897 = _T_234 ? _GEN_1882 : _GEN_1872; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 224:21]
  wire  _GEN_1898 = _T_371 | _GEN_1893; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 241:29]
  wire [63:0] _GEN_1899 = _T_371 ? _T_359 : _GEN_1894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 242:29]
  wire [63:0] _GEN_1900 = _T_371 ? _GEN_1895 : _T_359; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 244:26]
  wire  _GEN_1902 = _T_371 ? _GEN_1897 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 240:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1903 = $signed(_T_325) < $signed(_T_326) ? _GEN_1898 : _GEN_1893; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire [63:0] _GEN_1904 = $signed(_T_325) < $signed(_T_326) ? _GEN_1899 : _GEN_1894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire [63:0] _GEN_1905 = $signed(_T_325) < $signed(_T_326) ? _GEN_1900 : _GEN_1895; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire  _GEN_1907 = $signed(_T_325) < $signed(_T_326) ? _GEN_1902 : _GEN_1897; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 239:55]
  wire  _GEN_1918 = _T_261 ? _GEN_1903 : _GEN_1893; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire [63:0] _GEN_1919 = _T_261 ? _GEN_1904 : _GEN_1894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire [63:0] _GEN_1920 = _T_261 ? _GEN_1905 : _GEN_1895; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire  _GEN_1922 = _T_261 ? _GEN_1907 : _GEN_1897; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 237:21]
  wire  _GEN_1923 = _T_371 | _GEN_1918; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 253:29]
  wire [63:0] _GEN_1924 = _T_371 ? _T_359 : _GEN_1919; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 254:29]
  wire [63:0] _GEN_1925 = _T_371 ? _GEN_1920 : _T_359; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 256:26]
  wire  _GEN_1927 = _T_371 ? _GEN_1922 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 252:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1928 = _GEN_101 < _GEN_910 ? _GEN_1923 : _GEN_1918; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire [63:0] _GEN_1929 = _GEN_101 < _GEN_910 ? _GEN_1924 : _GEN_1919; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire [63:0] _GEN_1930 = _GEN_101 < _GEN_910 ? _GEN_1925 : _GEN_1920; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire  _GEN_1932 = _GEN_101 < _GEN_910 ? _GEN_1927 : _GEN_1922; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 251:41]
  wire  _GEN_1943 = _T_290 ? _GEN_1928 : _GEN_1918; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire [63:0] _GEN_1944 = _T_290 ? _GEN_1929 : _GEN_1919; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire [63:0] _GEN_1945 = _T_290 ? _GEN_1930 : _GEN_1920; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire  _GEN_1947 = _T_290 ? _GEN_1932 : _GEN_1922; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 249:22]
  wire  _GEN_1948 = _T_371 | _GEN_1943; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 266:29]
  wire [63:0] _GEN_1949 = _T_371 ? _T_359 : _GEN_1944; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 267:29]
  wire [63:0] _GEN_1950 = _T_371 ? _GEN_1945 : _T_359; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 269:26]
  wire  _GEN_1952 = _T_371 ? _GEN_1947 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 265:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1953 = $signed(_T_325) >= $signed(_T_326) ? _GEN_1948 : _GEN_1943; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire [63:0] _GEN_1954 = $signed(_T_325) >= $signed(_T_326) ? _GEN_1949 : _GEN_1944; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire [63:0] _GEN_1955 = $signed(_T_325) >= $signed(_T_326) ? _GEN_1950 : _GEN_1945; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire  _GEN_1957 = $signed(_T_325) >= $signed(_T_326) ? _GEN_1952 : _GEN_1947; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 264:56]
  wire  _GEN_1968 = _T_317 ? _GEN_1953 : _GEN_1943; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire [63:0] _GEN_1969 = _T_317 ? _GEN_1954 : _GEN_1944; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire [63:0] _GEN_1970 = _T_317 ? _GEN_1955 : _GEN_1945; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire  _GEN_1972 = _T_317 ? _GEN_1957 : _GEN_1947; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 262:21]
  wire  _GEN_1973 = _T_371 | _GEN_1968; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 278:29]
  wire [63:0] _GEN_1974 = _T_371 ? _T_359 : _GEN_1969; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 279:29]
  wire [63:0] _GEN_1975 = _T_371 ? _GEN_1970 : _T_359; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 281:26]
  wire  _GEN_1977 = _T_371 ? _GEN_1972 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 277:57 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_1978 = _GEN_101 >= _GEN_910 ? _GEN_1973 : _GEN_1968; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire [63:0] _GEN_1979 = _GEN_101 >= _GEN_910 ? _GEN_1974 : _GEN_1969; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire [63:0] _GEN_1980 = _GEN_101 >= _GEN_910 ? _GEN_1975 : _GEN_1970; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire  _GEN_1982 = _GEN_101 >= _GEN_910 ? _GEN_1977 : _GEN_1972; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 276:42]
  wire  _GEN_1993 = _T_346 ? _GEN_1978 : _GEN_1968; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire [63:0] _GEN_1994 = _T_346 ? _GEN_1979 : _GEN_1969; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire [63:0] _GEN_1995 = _T_346 ? _GEN_1980 : _GEN_1970; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire  _GEN_1997 = _T_346 ? _GEN_1982 : _GEN_1972; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 274:22]
  wire [5:0] next_reg_rOff = {_T_844[2:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 58:51]
  wire [63:0] next_reg_LevelVec__2_addr = {8'h0,io_now_csr_satp[43:0],_T_844[38:30],3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 268:31]
  wire [63:0] _next_reg_LevelVec_1_addr_T_3 = {8'h0,next_reg_PTE_30_ppn,_T_844[29:21],3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 302:54]
  wire [63:0] _GEN_1999 = next_reg_PTEFlag_30_r | next_reg_PTEFlag_30_x ? 64'h0 : _next_reg_LevelVec_1_addr_T_3; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 287:42 292:47 302:48]
  wire [63:0] next_reg_LevelVec__1_addr = ~next_reg_PTEFlag_30_v | ~next_reg_PTEFlag_30_r & next_reg_PTEFlag_30_w ? 64'h0
     : _GEN_1999; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 277:57 282:45]
  wire [63:0] _next_reg_LevelVec_0_addr_T_3 = {8'h0,next_reg_PTE_31_ppn,_T_844[20:12],3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 305:54]
  wire [63:0] _GEN_2014 = next_reg_PTEFlag_31_r | next_reg_PTEFlag_31_x ? 64'h0 : _next_reg_LevelVec_0_addr_T_3; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 287:42 292:47 305:48]
  wire [63:0] _GEN_2018 = ~next_reg_PTEFlag_31_v | ~next_reg_PTEFlag_31_r & next_reg_PTEFlag_31_w ? 64'h0 : _GEN_2014; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 277:57 282:45]
  wire [63:0] _GEN_2022 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec__1_addr : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] next_reg_LevelVec__0_addr = next_reg_LevelVec_10_1_valid ? _GEN_2018 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 271:41 317:43]
  wire [63:0] _GEN_2033 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec__0_addr : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [55:0] _next_reg_finaladdr_T_5 = {_GEN_8145[53:10],_T_844[11:0]}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 364:31]
  wire [43:0] _next_reg_finaladdr_T_6 = ~next_reg_mask_10; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 364:106]
  wire [55:0] _GEN_11189 = {{12'd0}, _next_reg_finaladdr_T_6}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 364:103]
  wire [55:0] _next_reg_finaladdr_T_7 = _next_reg_finaladdr_T_5 & _GEN_11189; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 364:103]
  wire [63:0] _GEN_11190 = {{20'd0}, next_reg_mask_10}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 366:26]
  wire [63:0] _next_reg_finaladdr_T_8 = _T_844 & _GEN_11190; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 366:26]
  wire [63:0] _GEN_11191 = {{8'd0}, _next_reg_finaladdr_T_7}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 366:18]
  wire [63:0] _next_reg_finaladdr_T_9 = _GEN_11191 | _next_reg_finaladdr_T_8; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 366:18]
  wire [63:0] _GEN_2059 = _next_reg_T_797 ? 64'h0 : _next_reg_finaladdr_T_9; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 349:99 352:26 364:23]
  wire [63:0] _GEN_2065 = next_reg_permLoad_10 ? _GEN_2059 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 346:11 372:24]
  wire [63:0] next_reg_finaladdr = ~(next_reg_successLevel_10 == 2'h3) ? _GEN_2065 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 335:37 377:22]
  wire [63:0] _GEN_2091 = next_reg_success_10 ? next_reg_finaladdr : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 69:25 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire  _GEN_2093 = next_reg_success_10 ? _GEN_1997 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [63:0] _GEN_2095 = next_reg_vmEnable_10 ? next_reg_LevelVec__2_addr : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_2097 = next_reg_vmEnable_10 & next_reg_LevelVec_10_1_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_2098 = next_reg_vmEnable_10 ? _GEN_2022 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_2100 = next_reg_vmEnable_10 & next_reg_LevelVec_10_0_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_2101 = next_reg_vmEnable_10 ? _GEN_2033 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_2107 = next_reg_vmEnable_10 ? _GEN_2091 : _T_844; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22 74:23]
  wire  _GEN_2109 = next_reg_vmEnable_10 ? _GEN_2093 : _GEN_1997; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _next_reg_T_100 = io_mem_read_data >> next_reg_rOff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 77:22]
  wire [63:0] _next_reg_T_101 = _next_reg_T_100 & 64'hff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 77:31]
  wire  next_reg_signBit = _next_reg_T_101[7]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [55:0] _next_reg_T_104 = next_reg_signBit ? 56'hffffffffffffff : 56'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_105 = {_next_reg_T_104,_next_reg_T_101[7:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_2111 = 5'h1 == rd ? _next_reg_T_105 : _GEN_1814; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2112 = 5'h2 == rd ? _next_reg_T_105 : _GEN_1815; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2113 = 5'h3 == rd ? _next_reg_T_105 : _GEN_1816; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2114 = 5'h4 == rd ? _next_reg_T_105 : _GEN_1817; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2115 = 5'h5 == rd ? _next_reg_T_105 : _GEN_1818; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2116 = 5'h6 == rd ? _next_reg_T_105 : _GEN_1819; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2117 = 5'h7 == rd ? _next_reg_T_105 : _GEN_1820; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2118 = 5'h8 == rd ? _next_reg_T_105 : _GEN_1821; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2119 = 5'h9 == rd ? _next_reg_T_105 : _GEN_1822; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2120 = 5'ha == rd ? _next_reg_T_105 : _GEN_1823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2121 = 5'hb == rd ? _next_reg_T_105 : _GEN_1824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2122 = 5'hc == rd ? _next_reg_T_105 : _GEN_1825; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2123 = 5'hd == rd ? _next_reg_T_105 : _GEN_1826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2124 = 5'he == rd ? _next_reg_T_105 : _GEN_1827; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2125 = 5'hf == rd ? _next_reg_T_105 : _GEN_1828; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2126 = 5'h10 == rd ? _next_reg_T_105 : _GEN_1829; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2127 = 5'h11 == rd ? _next_reg_T_105 : _GEN_1830; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2128 = 5'h12 == rd ? _next_reg_T_105 : _GEN_1831; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2129 = 5'h13 == rd ? _next_reg_T_105 : _GEN_1832; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2130 = 5'h14 == rd ? _next_reg_T_105 : _GEN_1833; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2131 = 5'h15 == rd ? _next_reg_T_105 : _GEN_1834; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2132 = 5'h16 == rd ? _next_reg_T_105 : _GEN_1835; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2133 = 5'h17 == rd ? _next_reg_T_105 : _GEN_1836; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2134 = 5'h18 == rd ? _next_reg_T_105 : _GEN_1837; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2135 = 5'h19 == rd ? _next_reg_T_105 : _GEN_1838; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2136 = 5'h1a == rd ? _next_reg_T_105 : _GEN_1839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2137 = 5'h1b == rd ? _next_reg_T_105 : _GEN_1840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2138 = 5'h1c == rd ? _next_reg_T_105 : _GEN_1841; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2139 = 5'h1d == rd ? _next_reg_T_105 : _GEN_1842; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2140 = 5'h1e == rd ? _next_reg_T_105 : _GEN_1843; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire [63:0] _GEN_2141 = 5'h1f == rd ? _next_reg_T_105 : _GEN_1844; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 291:{22,22}]
  wire  _GEN_2201 = _T_373 & next_reg_vmEnable_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2202 = _T_373 ? _GEN_2095 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire  _GEN_2204 = _T_373 & _GEN_2097; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2205 = _T_373 ? _GEN_2098 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire  _GEN_2207 = _T_373 & _GEN_2100; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2208 = _T_373 ? _GEN_2101 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2214 = _T_373 ? _GEN_2107 : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire  _GEN_2216 = _T_373 ? _GEN_2109 : _GEN_1997; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [6:0] _GEN_2217 = _T_373 ? 7'h8 : 7'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [63:0] _GEN_2219 = _T_373 ? _GEN_2111 : _GEN_1814; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2220 = _T_373 ? _GEN_2112 : _GEN_1815; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2221 = _T_373 ? _GEN_2113 : _GEN_1816; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2222 = _T_373 ? _GEN_2114 : _GEN_1817; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2223 = _T_373 ? _GEN_2115 : _GEN_1818; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2224 = _T_373 ? _GEN_2116 : _GEN_1819; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2225 = _T_373 ? _GEN_2117 : _GEN_1820; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2226 = _T_373 ? _GEN_2118 : _GEN_1821; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2227 = _T_373 ? _GEN_2119 : _GEN_1822; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2228 = _T_373 ? _GEN_2120 : _GEN_1823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2229 = _T_373 ? _GEN_2121 : _GEN_1824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2230 = _T_373 ? _GEN_2122 : _GEN_1825; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2231 = _T_373 ? _GEN_2123 : _GEN_1826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2232 = _T_373 ? _GEN_2124 : _GEN_1827; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2233 = _T_373 ? _GEN_2125 : _GEN_1828; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2234 = _T_373 ? _GEN_2126 : _GEN_1829; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2235 = _T_373 ? _GEN_2127 : _GEN_1830; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2236 = _T_373 ? _GEN_2128 : _GEN_1831; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2237 = _T_373 ? _GEN_2129 : _GEN_1832; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2238 = _T_373 ? _GEN_2130 : _GEN_1833; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2239 = _T_373 ? _GEN_2131 : _GEN_1834; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2240 = _T_373 ? _GEN_2132 : _GEN_1835; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2241 = _T_373 ? _GEN_2133 : _GEN_1836; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2242 = _T_373 ? _GEN_2134 : _GEN_1837; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2243 = _T_373 ? _GEN_2135 : _GEN_1838; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2244 = _T_373 ? _GEN_2136 : _GEN_1839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2245 = _T_373 ? _GEN_2137 : _GEN_1840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2246 = _T_373 ? _GEN_2138 : _GEN_1841; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2247 = _T_373 ? _GEN_2139 : _GEN_1842; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2248 = _T_373 ? _GEN_2140 : _GEN_1843; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire [63:0] _GEN_2249 = _T_373 ? _GEN_2141 : _GEN_1844; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 288:20]
  wire  _GEN_2274 = next_reg_LevelVec_10_1_valid | _GEN_2204; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_2275 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec__1_addr : _GEN_2205; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire  _GEN_2285 = next_reg_LevelVec_10_0_valid | _GEN_2207; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_2286 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec__0_addr : _GEN_2208; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] _GEN_2344 = next_reg_success_10 ? next_reg_finaladdr : _GEN_2214; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 69:25]
  wire  _GEN_2346 = next_reg_success_10 ? _GEN_2216 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_2347 = next_reg_vmEnable_10 | _GEN_2201; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_2348 = next_reg_vmEnable_10 ? next_reg_LevelVec__2_addr : _GEN_2202; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_2350 = next_reg_vmEnable_10 ? _GEN_2274 : _GEN_2204; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_2351 = next_reg_vmEnable_10 ? _GEN_2275 : _GEN_2205; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_2353 = next_reg_vmEnable_10 ? _GEN_2285 : _GEN_2207; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_2354 = next_reg_vmEnable_10 ? _GEN_2286 : _GEN_2208; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_2360 = next_reg_vmEnable_10 ? _GEN_2344 : _T_844; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22 74:23]
  wire  _GEN_2362 = next_reg_vmEnable_10 ? _GEN_2346 : _GEN_2216; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _next_reg_T_161 = _next_reg_T_100 & 64'hffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 77:31]
  wire  next_reg_signBit_1 = _next_reg_T_161[15]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [47:0] _next_reg_T_164 = next_reg_signBit_1 ? 48'hffffffffffff : 48'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_165 = {_next_reg_T_164,_next_reg_T_161[15:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_2364 = 5'h1 == rd ? _next_reg_T_165 : _GEN_2219; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2365 = 5'h2 == rd ? _next_reg_T_165 : _GEN_2220; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2366 = 5'h3 == rd ? _next_reg_T_165 : _GEN_2221; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2367 = 5'h4 == rd ? _next_reg_T_165 : _GEN_2222; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2368 = 5'h5 == rd ? _next_reg_T_165 : _GEN_2223; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2369 = 5'h6 == rd ? _next_reg_T_165 : _GEN_2224; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2370 = 5'h7 == rd ? _next_reg_T_165 : _GEN_2225; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2371 = 5'h8 == rd ? _next_reg_T_165 : _GEN_2226; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2372 = 5'h9 == rd ? _next_reg_T_165 : _GEN_2227; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2373 = 5'ha == rd ? _next_reg_T_165 : _GEN_2228; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2374 = 5'hb == rd ? _next_reg_T_165 : _GEN_2229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2375 = 5'hc == rd ? _next_reg_T_165 : _GEN_2230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2376 = 5'hd == rd ? _next_reg_T_165 : _GEN_2231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2377 = 5'he == rd ? _next_reg_T_165 : _GEN_2232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2378 = 5'hf == rd ? _next_reg_T_165 : _GEN_2233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2379 = 5'h10 == rd ? _next_reg_T_165 : _GEN_2234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2380 = 5'h11 == rd ? _next_reg_T_165 : _GEN_2235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2381 = 5'h12 == rd ? _next_reg_T_165 : _GEN_2236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2382 = 5'h13 == rd ? _next_reg_T_165 : _GEN_2237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2383 = 5'h14 == rd ? _next_reg_T_165 : _GEN_2238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2384 = 5'h15 == rd ? _next_reg_T_165 : _GEN_2239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2385 = 5'h16 == rd ? _next_reg_T_165 : _GEN_2240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2386 = 5'h17 == rd ? _next_reg_T_165 : _GEN_2241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2387 = 5'h18 == rd ? _next_reg_T_165 : _GEN_2242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2388 = 5'h19 == rd ? _next_reg_T_165 : _GEN_2243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2389 = 5'h1a == rd ? _next_reg_T_165 : _GEN_2244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2390 = 5'h1b == rd ? _next_reg_T_165 : _GEN_2245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2391 = 5'h1c == rd ? _next_reg_T_165 : _GEN_2246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2392 = 5'h1d == rd ? _next_reg_T_165 : _GEN_2247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2393 = 5'h1e == rd ? _next_reg_T_165 : _GEN_2248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire [63:0] _GEN_2394 = 5'h1f == rd ? _next_reg_T_165 : _GEN_2249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 301:{22,22}]
  wire  _GEN_2395 = _T_846 | _T_373; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 63:22]
  wire  _GEN_2396 = _T_846 ? _GEN_2347 : _GEN_2201; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2397 = _T_846 ? _GEN_2348 : _GEN_2202; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire  _GEN_2399 = _T_846 ? _GEN_2350 : _GEN_2204; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2400 = _T_846 ? _GEN_2351 : _GEN_2205; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire  _GEN_2402 = _T_846 ? _GEN_2353 : _GEN_2207; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2403 = _T_846 ? _GEN_2354 : _GEN_2208; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2409 = _T_846 ? _GEN_2360 : _T_844; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 303:23]
  wire  _GEN_2411 = _T_846 ? _GEN_2362 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [6:0] _GEN_2412 = _T_846 ? 7'h10 : _GEN_2217; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 76:25]
  wire [63:0] _GEN_2414 = _T_846 ? _GEN_2364 : _GEN_2219; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2415 = _T_846 ? _GEN_2365 : _GEN_2220; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2416 = _T_846 ? _GEN_2366 : _GEN_2221; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2417 = _T_846 ? _GEN_2367 : _GEN_2222; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2418 = _T_846 ? _GEN_2368 : _GEN_2223; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2419 = _T_846 ? _GEN_2369 : _GEN_2224; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2420 = _T_846 ? _GEN_2370 : _GEN_2225; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2421 = _T_846 ? _GEN_2371 : _GEN_2226; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2422 = _T_846 ? _GEN_2372 : _GEN_2227; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2423 = _T_846 ? _GEN_2373 : _GEN_2228; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2424 = _T_846 ? _GEN_2374 : _GEN_2229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2425 = _T_846 ? _GEN_2375 : _GEN_2230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2426 = _T_846 ? _GEN_2376 : _GEN_2231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2427 = _T_846 ? _GEN_2377 : _GEN_2232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2428 = _T_846 ? _GEN_2378 : _GEN_2233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2429 = _T_846 ? _GEN_2379 : _GEN_2234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2430 = _T_846 ? _GEN_2380 : _GEN_2235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2431 = _T_846 ? _GEN_2381 : _GEN_2236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2432 = _T_846 ? _GEN_2382 : _GEN_2237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2433 = _T_846 ? _GEN_2383 : _GEN_2238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2434 = _T_846 ? _GEN_2384 : _GEN_2239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2435 = _T_846 ? _GEN_2385 : _GEN_2240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2436 = _T_846 ? _GEN_2386 : _GEN_2241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2437 = _T_846 ? _GEN_2387 : _GEN_2242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2438 = _T_846 ? _GEN_2388 : _GEN_2243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2439 = _T_846 ? _GEN_2389 : _GEN_2244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2440 = _T_846 ? _GEN_2390 : _GEN_2245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2441 = _T_846 ? _GEN_2391 : _GEN_2246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2442 = _T_846 ? _GEN_2392 : _GEN_2247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2443 = _T_846 ? _GEN_2393 : _GEN_2248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire [63:0] _GEN_2444 = _T_846 ? _GEN_2394 : _GEN_2249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 300:55]
  wire  _GEN_2453 = _T_393 ? _GEN_2395 : _T_373; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire  _GEN_2454 = _T_393 ? _GEN_2396 : _GEN_2201; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2455 = _T_393 ? _GEN_2397 : _GEN_2202; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire  _GEN_2457 = _T_393 ? _GEN_2399 : _GEN_2204; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2458 = _T_393 ? _GEN_2400 : _GEN_2205; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire  _GEN_2460 = _T_393 ? _GEN_2402 : _GEN_2207; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2461 = _T_393 ? _GEN_2403 : _GEN_2208; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2467 = _T_393 ? _GEN_2409 : _GEN_2214; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire  _GEN_2469 = _T_393 ? _GEN_2411 : _GEN_2216; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [6:0] _GEN_2470 = _T_393 ? _GEN_2412 : _GEN_2217; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2472 = _T_393 ? _GEN_2414 : _GEN_2219; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2473 = _T_393 ? _GEN_2415 : _GEN_2220; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2474 = _T_393 ? _GEN_2416 : _GEN_2221; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2475 = _T_393 ? _GEN_2417 : _GEN_2222; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2476 = _T_393 ? _GEN_2418 : _GEN_2223; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2477 = _T_393 ? _GEN_2419 : _GEN_2224; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2478 = _T_393 ? _GEN_2420 : _GEN_2225; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2479 = _T_393 ? _GEN_2421 : _GEN_2226; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2480 = _T_393 ? _GEN_2422 : _GEN_2227; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2481 = _T_393 ? _GEN_2423 : _GEN_2228; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2482 = _T_393 ? _GEN_2424 : _GEN_2229; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2483 = _T_393 ? _GEN_2425 : _GEN_2230; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2484 = _T_393 ? _GEN_2426 : _GEN_2231; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2485 = _T_393 ? _GEN_2427 : _GEN_2232; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2486 = _T_393 ? _GEN_2428 : _GEN_2233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2487 = _T_393 ? _GEN_2429 : _GEN_2234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2488 = _T_393 ? _GEN_2430 : _GEN_2235; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2489 = _T_393 ? _GEN_2431 : _GEN_2236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2490 = _T_393 ? _GEN_2432 : _GEN_2237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2491 = _T_393 ? _GEN_2433 : _GEN_2238; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2492 = _T_393 ? _GEN_2434 : _GEN_2239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2493 = _T_393 ? _GEN_2435 : _GEN_2240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2494 = _T_393 ? _GEN_2436 : _GEN_2241; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2495 = _T_393 ? _GEN_2437 : _GEN_2242; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2496 = _T_393 ? _GEN_2438 : _GEN_2243; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2497 = _T_393 ? _GEN_2439 : _GEN_2244; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2498 = _T_393 ? _GEN_2440 : _GEN_2245; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2499 = _T_393 ? _GEN_2441 : _GEN_2246; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2500 = _T_393 ? _GEN_2442 : _GEN_2247; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2501 = _T_393 ? _GEN_2443 : _GEN_2248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire [63:0] _GEN_2502 = _T_393 ? _GEN_2444 : _GEN_2249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 298:20]
  wire  _GEN_2527 = next_reg_LevelVec_10_1_valid | _GEN_2457; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_2528 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec__1_addr : _GEN_2458; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire  _GEN_2538 = next_reg_LevelVec_10_0_valid | _GEN_2460; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_2539 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec__0_addr : _GEN_2461; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] _GEN_2597 = next_reg_success_10 ? next_reg_finaladdr : _GEN_2467; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 69:25]
  wire  _GEN_2599 = next_reg_success_10 ? _GEN_2469 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_2600 = next_reg_vmEnable_10 | _GEN_2454; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_2601 = next_reg_vmEnable_10 ? next_reg_LevelVec__2_addr : _GEN_2455; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_2603 = next_reg_vmEnable_10 ? _GEN_2527 : _GEN_2457; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_2604 = next_reg_vmEnable_10 ? _GEN_2528 : _GEN_2458; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_2606 = next_reg_vmEnable_10 ? _GEN_2538 : _GEN_2460; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_2607 = next_reg_vmEnable_10 ? _GEN_2539 : _GEN_2461; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_2613 = next_reg_vmEnable_10 ? _GEN_2597 : _T_844; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22 74:23]
  wire  _GEN_2615 = next_reg_vmEnable_10 ? _GEN_2599 : _GEN_2469; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _next_reg_T_221 = _next_reg_T_100 & 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 77:31]
  wire  next_reg_signBit_2 = _next_reg_T_221[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_224 = next_reg_signBit_2 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_225 = {_next_reg_T_224,_next_reg_T_221[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_2617 = 5'h1 == rd ? _next_reg_T_225 : _GEN_2472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2618 = 5'h2 == rd ? _next_reg_T_225 : _GEN_2473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2619 = 5'h3 == rd ? _next_reg_T_225 : _GEN_2474; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2620 = 5'h4 == rd ? _next_reg_T_225 : _GEN_2475; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2621 = 5'h5 == rd ? _next_reg_T_225 : _GEN_2476; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2622 = 5'h6 == rd ? _next_reg_T_225 : _GEN_2477; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2623 = 5'h7 == rd ? _next_reg_T_225 : _GEN_2478; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2624 = 5'h8 == rd ? _next_reg_T_225 : _GEN_2479; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2625 = 5'h9 == rd ? _next_reg_T_225 : _GEN_2480; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2626 = 5'ha == rd ? _next_reg_T_225 : _GEN_2481; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2627 = 5'hb == rd ? _next_reg_T_225 : _GEN_2482; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2628 = 5'hc == rd ? _next_reg_T_225 : _GEN_2483; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2629 = 5'hd == rd ? _next_reg_T_225 : _GEN_2484; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2630 = 5'he == rd ? _next_reg_T_225 : _GEN_2485; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2631 = 5'hf == rd ? _next_reg_T_225 : _GEN_2486; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2632 = 5'h10 == rd ? _next_reg_T_225 : _GEN_2487; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2633 = 5'h11 == rd ? _next_reg_T_225 : _GEN_2488; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2634 = 5'h12 == rd ? _next_reg_T_225 : _GEN_2489; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2635 = 5'h13 == rd ? _next_reg_T_225 : _GEN_2490; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2636 = 5'h14 == rd ? _next_reg_T_225 : _GEN_2491; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2637 = 5'h15 == rd ? _next_reg_T_225 : _GEN_2492; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2638 = 5'h16 == rd ? _next_reg_T_225 : _GEN_2493; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2639 = 5'h17 == rd ? _next_reg_T_225 : _GEN_2494; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2640 = 5'h18 == rd ? _next_reg_T_225 : _GEN_2495; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2641 = 5'h19 == rd ? _next_reg_T_225 : _GEN_2496; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2642 = 5'h1a == rd ? _next_reg_T_225 : _GEN_2497; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2643 = 5'h1b == rd ? _next_reg_T_225 : _GEN_2498; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2644 = 5'h1c == rd ? _next_reg_T_225 : _GEN_2499; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2645 = 5'h1d == rd ? _next_reg_T_225 : _GEN_2500; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2646 = 5'h1e == rd ? _next_reg_T_225 : _GEN_2501; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire [63:0] _GEN_2647 = 5'h1f == rd ? _next_reg_T_225 : _GEN_2502; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 310:{22,22}]
  wire  _GEN_2648 = _T_848 | _GEN_2453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 63:22]
  wire  _GEN_2649 = _T_848 ? _GEN_2600 : _GEN_2454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2650 = _T_848 ? _GEN_2601 : _GEN_2455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire  _GEN_2652 = _T_848 ? _GEN_2603 : _GEN_2457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2653 = _T_848 ? _GEN_2604 : _GEN_2458; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire  _GEN_2655 = _T_848 ? _GEN_2606 : _GEN_2460; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2656 = _T_848 ? _GEN_2607 : _GEN_2461; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2662 = _T_848 ? _GEN_2613 : _T_844; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 312:23]
  wire  _GEN_2664 = _T_848 ? _GEN_2615 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [6:0] _GEN_2665 = _T_848 ? 7'h20 : _GEN_2470; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 76:25]
  wire [63:0] _GEN_2667 = _T_848 ? _GEN_2617 : _GEN_2472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2668 = _T_848 ? _GEN_2618 : _GEN_2473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2669 = _T_848 ? _GEN_2619 : _GEN_2474; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2670 = _T_848 ? _GEN_2620 : _GEN_2475; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2671 = _T_848 ? _GEN_2621 : _GEN_2476; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2672 = _T_848 ? _GEN_2622 : _GEN_2477; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2673 = _T_848 ? _GEN_2623 : _GEN_2478; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2674 = _T_848 ? _GEN_2624 : _GEN_2479; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2675 = _T_848 ? _GEN_2625 : _GEN_2480; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2676 = _T_848 ? _GEN_2626 : _GEN_2481; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2677 = _T_848 ? _GEN_2627 : _GEN_2482; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2678 = _T_848 ? _GEN_2628 : _GEN_2483; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2679 = _T_848 ? _GEN_2629 : _GEN_2484; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2680 = _T_848 ? _GEN_2630 : _GEN_2485; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2681 = _T_848 ? _GEN_2631 : _GEN_2486; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2682 = _T_848 ? _GEN_2632 : _GEN_2487; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2683 = _T_848 ? _GEN_2633 : _GEN_2488; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2684 = _T_848 ? _GEN_2634 : _GEN_2489; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2685 = _T_848 ? _GEN_2635 : _GEN_2490; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2686 = _T_848 ? _GEN_2636 : _GEN_2491; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2687 = _T_848 ? _GEN_2637 : _GEN_2492; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2688 = _T_848 ? _GEN_2638 : _GEN_2493; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2689 = _T_848 ? _GEN_2639 : _GEN_2494; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2690 = _T_848 ? _GEN_2640 : _GEN_2495; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2691 = _T_848 ? _GEN_2641 : _GEN_2496; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2692 = _T_848 ? _GEN_2642 : _GEN_2497; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2693 = _T_848 ? _GEN_2643 : _GEN_2498; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2694 = _T_848 ? _GEN_2644 : _GEN_2499; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2695 = _T_848 ? _GEN_2645 : _GEN_2500; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2696 = _T_848 ? _GEN_2646 : _GEN_2501; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire [63:0] _GEN_2697 = _T_848 ? _GEN_2647 : _GEN_2502; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 309:55]
  wire  _GEN_2706 = _T_413 ? _GEN_2648 : _GEN_2453; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2707 = _T_413 ? _GEN_2649 : _GEN_2454; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2708 = _T_413 ? _GEN_2650 : _GEN_2455; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2710 = _T_413 ? _GEN_2652 : _GEN_2457; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2711 = _T_413 ? _GEN_2653 : _GEN_2458; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2713 = _T_413 ? _GEN_2655 : _GEN_2460; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2714 = _T_413 ? _GEN_2656 : _GEN_2461; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2720 = _T_413 ? _GEN_2662 : _GEN_2467; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2722 = _T_413 ? _GEN_2664 : _GEN_2469; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [6:0] _GEN_2723 = _T_413 ? _GEN_2665 : _GEN_2470; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2725 = _T_413 ? _GEN_2667 : _GEN_2472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2726 = _T_413 ? _GEN_2668 : _GEN_2473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2727 = _T_413 ? _GEN_2669 : _GEN_2474; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2728 = _T_413 ? _GEN_2670 : _GEN_2475; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2729 = _T_413 ? _GEN_2671 : _GEN_2476; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2730 = _T_413 ? _GEN_2672 : _GEN_2477; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2731 = _T_413 ? _GEN_2673 : _GEN_2478; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2732 = _T_413 ? _GEN_2674 : _GEN_2479; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2733 = _T_413 ? _GEN_2675 : _GEN_2480; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2734 = _T_413 ? _GEN_2676 : _GEN_2481; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2735 = _T_413 ? _GEN_2677 : _GEN_2482; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2736 = _T_413 ? _GEN_2678 : _GEN_2483; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2737 = _T_413 ? _GEN_2679 : _GEN_2484; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2738 = _T_413 ? _GEN_2680 : _GEN_2485; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2739 = _T_413 ? _GEN_2681 : _GEN_2486; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2740 = _T_413 ? _GEN_2682 : _GEN_2487; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2741 = _T_413 ? _GEN_2683 : _GEN_2488; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2742 = _T_413 ? _GEN_2684 : _GEN_2489; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2743 = _T_413 ? _GEN_2685 : _GEN_2490; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2744 = _T_413 ? _GEN_2686 : _GEN_2491; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2745 = _T_413 ? _GEN_2687 : _GEN_2492; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2746 = _T_413 ? _GEN_2688 : _GEN_2493; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2747 = _T_413 ? _GEN_2689 : _GEN_2494; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2748 = _T_413 ? _GEN_2690 : _GEN_2495; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2749 = _T_413 ? _GEN_2691 : _GEN_2496; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2750 = _T_413 ? _GEN_2692 : _GEN_2497; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2751 = _T_413 ? _GEN_2693 : _GEN_2498; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2752 = _T_413 ? _GEN_2694 : _GEN_2499; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2753 = _T_413 ? _GEN_2695 : _GEN_2500; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2754 = _T_413 ? _GEN_2696 : _GEN_2501; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire [63:0] _GEN_2755 = _T_413 ? _GEN_2697 : _GEN_2502; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 307:20]
  wire  _GEN_2782 = next_reg_LevelVec_10_1_valid | _GEN_2710; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_2783 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec__1_addr : _GEN_2711; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire  _GEN_2793 = next_reg_LevelVec_10_0_valid | _GEN_2713; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_2794 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec__0_addr : _GEN_2714; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] _GEN_2852 = next_reg_success_10 ? next_reg_finaladdr : _GEN_2720; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 69:25]
  wire  _GEN_2854 = next_reg_success_10 ? _GEN_2722 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_2855 = next_reg_vmEnable_10 | _GEN_2707; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_2856 = next_reg_vmEnable_10 ? next_reg_LevelVec__2_addr : _GEN_2708; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_2858 = next_reg_vmEnable_10 ? _GEN_2782 : _GEN_2710; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_2859 = next_reg_vmEnable_10 ? _GEN_2783 : _GEN_2711; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_2861 = next_reg_vmEnable_10 ? _GEN_2793 : _GEN_2713; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_2862 = next_reg_vmEnable_10 ? _GEN_2794 : _GEN_2714; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_2868 = next_reg_vmEnable_10 ? _GEN_2852 : _T_844; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22 74:23]
  wire  _GEN_2870 = next_reg_vmEnable_10 ? _GEN_2854 : _GEN_2722; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _next_reg_T_283 = {56'h0,_next_reg_T_101[7:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [63:0] _GEN_2872 = 5'h1 == rd ? _next_reg_T_283 : _GEN_2725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2873 = 5'h2 == rd ? _next_reg_T_283 : _GEN_2726; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2874 = 5'h3 == rd ? _next_reg_T_283 : _GEN_2727; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2875 = 5'h4 == rd ? _next_reg_T_283 : _GEN_2728; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2876 = 5'h5 == rd ? _next_reg_T_283 : _GEN_2729; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2877 = 5'h6 == rd ? _next_reg_T_283 : _GEN_2730; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2878 = 5'h7 == rd ? _next_reg_T_283 : _GEN_2731; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2879 = 5'h8 == rd ? _next_reg_T_283 : _GEN_2732; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2880 = 5'h9 == rd ? _next_reg_T_283 : _GEN_2733; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2881 = 5'ha == rd ? _next_reg_T_283 : _GEN_2734; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2882 = 5'hb == rd ? _next_reg_T_283 : _GEN_2735; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2883 = 5'hc == rd ? _next_reg_T_283 : _GEN_2736; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2884 = 5'hd == rd ? _next_reg_T_283 : _GEN_2737; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2885 = 5'he == rd ? _next_reg_T_283 : _GEN_2738; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2886 = 5'hf == rd ? _next_reg_T_283 : _GEN_2739; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2887 = 5'h10 == rd ? _next_reg_T_283 : _GEN_2740; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2888 = 5'h11 == rd ? _next_reg_T_283 : _GEN_2741; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2889 = 5'h12 == rd ? _next_reg_T_283 : _GEN_2742; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2890 = 5'h13 == rd ? _next_reg_T_283 : _GEN_2743; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2891 = 5'h14 == rd ? _next_reg_T_283 : _GEN_2744; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2892 = 5'h15 == rd ? _next_reg_T_283 : _GEN_2745; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2893 = 5'h16 == rd ? _next_reg_T_283 : _GEN_2746; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2894 = 5'h17 == rd ? _next_reg_T_283 : _GEN_2747; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2895 = 5'h18 == rd ? _next_reg_T_283 : _GEN_2748; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2896 = 5'h19 == rd ? _next_reg_T_283 : _GEN_2749; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2897 = 5'h1a == rd ? _next_reg_T_283 : _GEN_2750; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2898 = 5'h1b == rd ? _next_reg_T_283 : _GEN_2751; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2899 = 5'h1c == rd ? _next_reg_T_283 : _GEN_2752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2900 = 5'h1d == rd ? _next_reg_T_283 : _GEN_2753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2901 = 5'h1e == rd ? _next_reg_T_283 : _GEN_2754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire [63:0] _GEN_2902 = 5'h1f == rd ? _next_reg_T_283 : _GEN_2755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:{86,86}]
  wire  _GEN_2911 = _T_433 ? _GEN_2870 : _GEN_2722; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire  _GEN_2912 = _T_433 | _GEN_2706; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/LoadStore.scala 63:22]
  wire  _GEN_2913 = _T_433 ? _GEN_2855 : _GEN_2707; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2914 = _T_433 ? _GEN_2856 : _GEN_2708; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire  _GEN_2916 = _T_433 ? _GEN_2858 : _GEN_2710; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2917 = _T_433 ? _GEN_2859 : _GEN_2711; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire  _GEN_2919 = _T_433 ? _GEN_2861 : _GEN_2713; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2920 = _T_433 ? _GEN_2862 : _GEN_2714; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2926 = _T_433 ? _GEN_2868 : _GEN_2720; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [6:0] _GEN_2928 = _T_433 ? 7'h8 : _GEN_2723; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21 src/main/scala/rvspeccore/core/tool/LoadStore.scala 76:25]
  wire [63:0] _GEN_2930 = _T_433 ? _GEN_2872 : _GEN_2725; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2931 = _T_433 ? _GEN_2873 : _GEN_2726; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2932 = _T_433 ? _GEN_2874 : _GEN_2727; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2933 = _T_433 ? _GEN_2875 : _GEN_2728; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2934 = _T_433 ? _GEN_2876 : _GEN_2729; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2935 = _T_433 ? _GEN_2877 : _GEN_2730; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2936 = _T_433 ? _GEN_2878 : _GEN_2731; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2937 = _T_433 ? _GEN_2879 : _GEN_2732; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2938 = _T_433 ? _GEN_2880 : _GEN_2733; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2939 = _T_433 ? _GEN_2881 : _GEN_2734; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2940 = _T_433 ? _GEN_2882 : _GEN_2735; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2941 = _T_433 ? _GEN_2883 : _GEN_2736; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2942 = _T_433 ? _GEN_2884 : _GEN_2737; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2943 = _T_433 ? _GEN_2885 : _GEN_2738; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2944 = _T_433 ? _GEN_2886 : _GEN_2739; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2945 = _T_433 ? _GEN_2887 : _GEN_2740; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2946 = _T_433 ? _GEN_2888 : _GEN_2741; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2947 = _T_433 ? _GEN_2889 : _GEN_2742; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2948 = _T_433 ? _GEN_2890 : _GEN_2743; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2949 = _T_433 ? _GEN_2891 : _GEN_2744; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2950 = _T_433 ? _GEN_2892 : _GEN_2745; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2951 = _T_433 ? _GEN_2893 : _GEN_2746; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2952 = _T_433 ? _GEN_2894 : _GEN_2747; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2953 = _T_433 ? _GEN_2895 : _GEN_2748; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2954 = _T_433 ? _GEN_2896 : _GEN_2749; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2955 = _T_433 ? _GEN_2897 : _GEN_2750; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2956 = _T_433 ? _GEN_2898 : _GEN_2751; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2957 = _T_433 ? _GEN_2899 : _GEN_2752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2958 = _T_433 ? _GEN_2900 : _GEN_2753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2959 = _T_433 ? _GEN_2901 : _GEN_2754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire [63:0] _GEN_2960 = _T_433 ? _GEN_2902 : _GEN_2755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 316:21]
  wire  _GEN_2984 = next_reg_LevelVec_10_1_valid | _GEN_2916; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_2985 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec__1_addr : _GEN_2917; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire  _GEN_2995 = next_reg_LevelVec_10_0_valid | _GEN_2919; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_2996 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec__0_addr : _GEN_2920; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] _GEN_3054 = next_reg_success_10 ? next_reg_finaladdr : _GEN_2926; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 69:25]
  wire  _GEN_3056 = next_reg_success_10 ? _GEN_2911 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_3057 = next_reg_vmEnable_10 | _GEN_2913; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_3058 = next_reg_vmEnable_10 ? next_reg_LevelVec__2_addr : _GEN_2914; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_3060 = next_reg_vmEnable_10 ? _GEN_2984 : _GEN_2916; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_3061 = next_reg_vmEnable_10 ? _GEN_2985 : _GEN_2917; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_3063 = next_reg_vmEnable_10 ? _GEN_2995 : _GEN_2919; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_3064 = next_reg_vmEnable_10 ? _GEN_2996 : _GEN_2920; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_3070 = next_reg_vmEnable_10 ? _GEN_3054 : _T_844; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22 74:23]
  wire  _GEN_3072 = next_reg_vmEnable_10 ? _GEN_3056 : _GEN_2911; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _next_reg_T_341 = {48'h0,_next_reg_T_161[15:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [63:0] _GEN_3074 = 5'h1 == rd ? _next_reg_T_341 : _GEN_2930; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3075 = 5'h2 == rd ? _next_reg_T_341 : _GEN_2931; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3076 = 5'h3 == rd ? _next_reg_T_341 : _GEN_2932; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3077 = 5'h4 == rd ? _next_reg_T_341 : _GEN_2933; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3078 = 5'h5 == rd ? _next_reg_T_341 : _GEN_2934; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3079 = 5'h6 == rd ? _next_reg_T_341 : _GEN_2935; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3080 = 5'h7 == rd ? _next_reg_T_341 : _GEN_2936; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3081 = 5'h8 == rd ? _next_reg_T_341 : _GEN_2937; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3082 = 5'h9 == rd ? _next_reg_T_341 : _GEN_2938; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3083 = 5'ha == rd ? _next_reg_T_341 : _GEN_2939; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3084 = 5'hb == rd ? _next_reg_T_341 : _GEN_2940; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3085 = 5'hc == rd ? _next_reg_T_341 : _GEN_2941; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3086 = 5'hd == rd ? _next_reg_T_341 : _GEN_2942; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3087 = 5'he == rd ? _next_reg_T_341 : _GEN_2943; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3088 = 5'hf == rd ? _next_reg_T_341 : _GEN_2944; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3089 = 5'h10 == rd ? _next_reg_T_341 : _GEN_2945; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3090 = 5'h11 == rd ? _next_reg_T_341 : _GEN_2946; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3091 = 5'h12 == rd ? _next_reg_T_341 : _GEN_2947; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3092 = 5'h13 == rd ? _next_reg_T_341 : _GEN_2948; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3093 = 5'h14 == rd ? _next_reg_T_341 : _GEN_2949; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3094 = 5'h15 == rd ? _next_reg_T_341 : _GEN_2950; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3095 = 5'h16 == rd ? _next_reg_T_341 : _GEN_2951; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3096 = 5'h17 == rd ? _next_reg_T_341 : _GEN_2952; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3097 = 5'h18 == rd ? _next_reg_T_341 : _GEN_2953; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3098 = 5'h19 == rd ? _next_reg_T_341 : _GEN_2954; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3099 = 5'h1a == rd ? _next_reg_T_341 : _GEN_2955; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3100 = 5'h1b == rd ? _next_reg_T_341 : _GEN_2956; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3101 = 5'h1c == rd ? _next_reg_T_341 : _GEN_2957; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3102 = 5'h1d == rd ? _next_reg_T_341 : _GEN_2958; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3103 = 5'h1e == rd ? _next_reg_T_341 : _GEN_2959; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire [63:0] _GEN_3104 = 5'h1f == rd ? _next_reg_T_341 : _GEN_2960; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 320:{22,22}]
  wire  _GEN_3105 = _T_846 | _GEN_2912; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 63:22]
  wire  _GEN_3106 = _T_846 ? _GEN_3057 : _GEN_2913; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3107 = _T_846 ? _GEN_3058 : _GEN_2914; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire  _GEN_3109 = _T_846 ? _GEN_3060 : _GEN_2916; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3110 = _T_846 ? _GEN_3061 : _GEN_2917; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire  _GEN_3112 = _T_846 ? _GEN_3063 : _GEN_2919; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3113 = _T_846 ? _GEN_3064 : _GEN_2920; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3119 = _T_846 ? _GEN_3070 : _T_844; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 322:23]
  wire  _GEN_3121 = _T_846 ? _GEN_3072 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [6:0] _GEN_3122 = _T_846 ? 7'h10 : _GEN_2928; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 76:25]
  wire [63:0] _GEN_3124 = _T_846 ? _GEN_3074 : _GEN_2930; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3125 = _T_846 ? _GEN_3075 : _GEN_2931; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3126 = _T_846 ? _GEN_3076 : _GEN_2932; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3127 = _T_846 ? _GEN_3077 : _GEN_2933; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3128 = _T_846 ? _GEN_3078 : _GEN_2934; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3129 = _T_846 ? _GEN_3079 : _GEN_2935; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3130 = _T_846 ? _GEN_3080 : _GEN_2936; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3131 = _T_846 ? _GEN_3081 : _GEN_2937; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3132 = _T_846 ? _GEN_3082 : _GEN_2938; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3133 = _T_846 ? _GEN_3083 : _GEN_2939; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3134 = _T_846 ? _GEN_3084 : _GEN_2940; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3135 = _T_846 ? _GEN_3085 : _GEN_2941; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3136 = _T_846 ? _GEN_3086 : _GEN_2942; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3137 = _T_846 ? _GEN_3087 : _GEN_2943; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3138 = _T_846 ? _GEN_3088 : _GEN_2944; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3139 = _T_846 ? _GEN_3089 : _GEN_2945; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3140 = _T_846 ? _GEN_3090 : _GEN_2946; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3141 = _T_846 ? _GEN_3091 : _GEN_2947; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3142 = _T_846 ? _GEN_3092 : _GEN_2948; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3143 = _T_846 ? _GEN_3093 : _GEN_2949; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3144 = _T_846 ? _GEN_3094 : _GEN_2950; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3145 = _T_846 ? _GEN_3095 : _GEN_2951; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3146 = _T_846 ? _GEN_3096 : _GEN_2952; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3147 = _T_846 ? _GEN_3097 : _GEN_2953; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3148 = _T_846 ? _GEN_3098 : _GEN_2954; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3149 = _T_846 ? _GEN_3099 : _GEN_2955; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3150 = _T_846 ? _GEN_3100 : _GEN_2956; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3151 = _T_846 ? _GEN_3101 : _GEN_2957; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3152 = _T_846 ? _GEN_3102 : _GEN_2958; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3153 = _T_846 ? _GEN_3103 : _GEN_2959; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire [63:0] _GEN_3154 = _T_846 ? _GEN_3104 : _GEN_2960; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 319:55]
  wire  _GEN_3163 = _T_452 ? _GEN_3105 : _GEN_2912; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire  _GEN_3164 = _T_452 ? _GEN_3106 : _GEN_2913; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3165 = _T_452 ? _GEN_3107 : _GEN_2914; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire  _GEN_3167 = _T_452 ? _GEN_3109 : _GEN_2916; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3168 = _T_452 ? _GEN_3110 : _GEN_2917; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire  _GEN_3170 = _T_452 ? _GEN_3112 : _GEN_2919; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3171 = _T_452 ? _GEN_3113 : _GEN_2920; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3177 = _T_452 ? _GEN_3119 : _GEN_2926; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire  _GEN_3179 = _T_452 ? _GEN_3121 : _GEN_2911; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [6:0] _GEN_3180 = _T_452 ? _GEN_3122 : _GEN_2928; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3182 = _T_452 ? _GEN_3124 : _GEN_2930; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3183 = _T_452 ? _GEN_3125 : _GEN_2931; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3184 = _T_452 ? _GEN_3126 : _GEN_2932; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3185 = _T_452 ? _GEN_3127 : _GEN_2933; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3186 = _T_452 ? _GEN_3128 : _GEN_2934; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3187 = _T_452 ? _GEN_3129 : _GEN_2935; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3188 = _T_452 ? _GEN_3130 : _GEN_2936; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3189 = _T_452 ? _GEN_3131 : _GEN_2937; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3190 = _T_452 ? _GEN_3132 : _GEN_2938; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3191 = _T_452 ? _GEN_3133 : _GEN_2939; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3192 = _T_452 ? _GEN_3134 : _GEN_2940; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3193 = _T_452 ? _GEN_3135 : _GEN_2941; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3194 = _T_452 ? _GEN_3136 : _GEN_2942; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3195 = _T_452 ? _GEN_3137 : _GEN_2943; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3196 = _T_452 ? _GEN_3138 : _GEN_2944; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3197 = _T_452 ? _GEN_3139 : _GEN_2945; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3198 = _T_452 ? _GEN_3140 : _GEN_2946; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3199 = _T_452 ? _GEN_3141 : _GEN_2947; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3200 = _T_452 ? _GEN_3142 : _GEN_2948; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3201 = _T_452 ? _GEN_3143 : _GEN_2949; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3202 = _T_452 ? _GEN_3144 : _GEN_2950; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3203 = _T_452 ? _GEN_3145 : _GEN_2951; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3204 = _T_452 ? _GEN_3146 : _GEN_2952; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3205 = _T_452 ? _GEN_3147 : _GEN_2953; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3206 = _T_452 ? _GEN_3148 : _GEN_2954; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3207 = _T_452 ? _GEN_3149 : _GEN_2955; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3208 = _T_452 ? _GEN_3150 : _GEN_2956; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3209 = _T_452 ? _GEN_3151 : _GEN_2957; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3210 = _T_452 ? _GEN_3152 : _GEN_2958; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3211 = _T_452 ? _GEN_3153 : _GEN_2959; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire [63:0] _GEN_3212 = _T_452 ? _GEN_3154 : _GEN_2960; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 317:21]
  wire  _GEN_3239 = next_reg_LevelVec_10_1_valid | _GEN_3167; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_3240 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec__1_addr : _GEN_3168; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire  _GEN_3250 = next_reg_LevelVec_10_0_valid | _GEN_3170; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_3251 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec__0_addr : _GEN_3171; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] _GEN_3283 = next_reg_permStore_10 ? _GEN_2059 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 346:11 372:24]
  wire [63:0] finaladdr_1 = ~(next_reg_successLevel_10 == 2'h3) ? _GEN_3283 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 335:37 377:22]
  wire [63:0] _GEN_3309 = success_8 ? finaladdr_1 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 97:26 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire  _GEN_3311 = success_8 ? _GEN_3179 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_3312 = next_reg_vmEnable_10 | _GEN_3164; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_3313 = next_reg_vmEnable_10 ? next_reg_LevelVec__2_addr : _GEN_3165; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_3315 = next_reg_vmEnable_10 ? _GEN_3239 : _GEN_3167; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_3316 = next_reg_vmEnable_10 ? _GEN_3240 : _GEN_3168; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_3318 = next_reg_vmEnable_10 ? _GEN_3250 : _GEN_3170; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_3319 = next_reg_vmEnable_10 ? _GEN_3251 : _GEN_3171; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_3325 = next_reg_vmEnable_10 ? _GEN_3309 : _T_844; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22 102:24]
  wire  _GEN_3327 = next_reg_vmEnable_10 ? _GEN_3311 : _GEN_3179; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_3337 = _T_472 ? _GEN_3327 : _GEN_3179; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20]
  wire  _GEN_3339 = _T_472 ? _GEN_3312 : _GEN_3164; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20]
  wire [63:0] _GEN_3340 = _T_472 ? _GEN_3313 : _GEN_3165; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20]
  wire  _GEN_3342 = _T_472 ? _GEN_3315 : _GEN_3167; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20]
  wire [63:0] _GEN_3343 = _T_472 ? _GEN_3316 : _GEN_3168; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20]
  wire  _GEN_3345 = _T_472 ? _GEN_3318 : _GEN_3170; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20]
  wire [63:0] _GEN_3346 = _T_472 ? _GEN_3319 : _GEN_3171; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20]
  wire [63:0] _GEN_3352 = _T_472 ? _GEN_3325 : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [6:0] _GEN_3354 = _T_472 ? 7'h8 : 7'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/LoadStore.scala 104:26 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire [63:0] _GEN_3355 = _T_472 ? {{56'd0}, _GEN_910[7:0]} : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 327:20 src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:26 src/main/scala/rvspeccore/core/RiscvCore.scala 119:7]
  wire  _GEN_3379 = next_reg_LevelVec_10_1_valid | _GEN_3342; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_3380 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec__1_addr : _GEN_3343; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire  _GEN_3390 = next_reg_LevelVec_10_0_valid | _GEN_3345; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_3391 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec__0_addr : _GEN_3346; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] _GEN_3449 = success_8 ? finaladdr_1 : _GEN_3352; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 97:26]
  wire  _GEN_3451 = success_8 ? _GEN_3337 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_3452 = next_reg_vmEnable_10 | _GEN_3339; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_3453 = next_reg_vmEnable_10 ? next_reg_LevelVec__2_addr : _GEN_3340; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_3455 = next_reg_vmEnable_10 ? _GEN_3379 : _GEN_3342; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_3456 = next_reg_vmEnable_10 ? _GEN_3380 : _GEN_3343; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_3458 = next_reg_vmEnable_10 ? _GEN_3390 : _GEN_3345; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_3459 = next_reg_vmEnable_10 ? _GEN_3391 : _GEN_3346; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_3465 = next_reg_vmEnable_10 ? _GEN_3449 : _T_844; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22 102:24]
  wire  _GEN_3467 = next_reg_vmEnable_10 ? _GEN_3451 : _GEN_3337; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_3468 = _T_846 | _T_472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 92:23]
  wire  _GEN_3469 = _T_846 ? _GEN_3452 : _GEN_3339; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55]
  wire [63:0] _GEN_3470 = _T_846 ? _GEN_3453 : _GEN_3340; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55]
  wire  _GEN_3472 = _T_846 ? _GEN_3455 : _GEN_3342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55]
  wire [63:0] _GEN_3473 = _T_846 ? _GEN_3456 : _GEN_3343; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55]
  wire  _GEN_3475 = _T_846 ? _GEN_3458 : _GEN_3345; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55]
  wire [63:0] _GEN_3476 = _T_846 ? _GEN_3459 : _GEN_3346; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55]
  wire [63:0] _GEN_3482 = _T_846 ? _GEN_3465 : _T_844; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 333:24]
  wire  _GEN_3484 = _T_846 ? _GEN_3467 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [6:0] _GEN_3485 = _T_846 ? 7'h10 : _GEN_3354; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 104:26]
  wire [63:0] _GEN_3486 = _T_846 ? {{48'd0}, _GEN_910[15:0]} : _GEN_3355; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 330:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:26]
  wire  _GEN_3496 = _T_547 ? _GEN_3468 : _T_472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire  _GEN_3497 = _T_547 ? _GEN_3469 : _GEN_3339; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [63:0] _GEN_3498 = _T_547 ? _GEN_3470 : _GEN_3340; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire  _GEN_3500 = _T_547 ? _GEN_3472 : _GEN_3342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [63:0] _GEN_3501 = _T_547 ? _GEN_3473 : _GEN_3343; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire  _GEN_3503 = _T_547 ? _GEN_3475 : _GEN_3345; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [63:0] _GEN_3504 = _T_547 ? _GEN_3476 : _GEN_3346; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [63:0] _GEN_3510 = _T_547 ? _GEN_3482 : _GEN_3352; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire  _GEN_3512 = _T_547 ? _GEN_3484 : _GEN_3337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [6:0] _GEN_3513 = _T_547 ? _GEN_3485 : _GEN_3354; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire [63:0] _GEN_3514 = _T_547 ? _GEN_3486 : _GEN_3355; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 328:20]
  wire  _GEN_3539 = next_reg_LevelVec_10_1_valid | _GEN_3500; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_3540 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec__1_addr : _GEN_3501; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire  _GEN_3550 = next_reg_LevelVec_10_0_valid | _GEN_3503; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_3551 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec__0_addr : _GEN_3504; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] _GEN_3609 = success_8 ? finaladdr_1 : _GEN_3510; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 97:26]
  wire  _GEN_3611 = success_8 ? _GEN_3512 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_3612 = next_reg_vmEnable_10 | _GEN_3497; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_3613 = next_reg_vmEnable_10 ? next_reg_LevelVec__2_addr : _GEN_3498; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_3615 = next_reg_vmEnable_10 ? _GEN_3539 : _GEN_3500; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_3616 = next_reg_vmEnable_10 ? _GEN_3540 : _GEN_3501; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_3618 = next_reg_vmEnable_10 ? _GEN_3550 : _GEN_3503; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_3619 = next_reg_vmEnable_10 ? _GEN_3551 : _GEN_3504; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_3625 = next_reg_vmEnable_10 ? _GEN_3609 : _T_844; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22 102:24]
  wire  _GEN_3627 = next_reg_vmEnable_10 ? _GEN_3611 : _GEN_3512; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_3628 = _T_848 | _GEN_3496; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 92:23]
  wire  _GEN_3629 = _T_848 ? _GEN_3612 : _GEN_3497; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55]
  wire [63:0] _GEN_3630 = _T_848 ? _GEN_3613 : _GEN_3498; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55]
  wire  _GEN_3632 = _T_848 ? _GEN_3615 : _GEN_3500; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55]
  wire [63:0] _GEN_3633 = _T_848 ? _GEN_3616 : _GEN_3501; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55]
  wire  _GEN_3635 = _T_848 ? _GEN_3618 : _GEN_3503; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55]
  wire [63:0] _GEN_3636 = _T_848 ? _GEN_3619 : _GEN_3504; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55]
  wire [63:0] _GEN_3642 = _T_848 ? _GEN_3625 : _T_844; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 342:24]
  wire  _GEN_3644 = _T_848 ? _GEN_3627 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [6:0] _GEN_3645 = _T_848 ? 7'h20 : _GEN_3513; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 104:26]
  wire [63:0] _GEN_3646 = _T_848 ? {{32'd0}, _GEN_910[31:0]} : _GEN_3514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 339:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:26]
  wire  _GEN_3656 = _T_623 ? _GEN_3628 : _GEN_3496; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire  _GEN_3657 = _T_623 ? _GEN_3629 : _GEN_3497; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [63:0] _GEN_3658 = _T_623 ? _GEN_3630 : _GEN_3498; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire  _GEN_3660 = _T_623 ? _GEN_3632 : _GEN_3500; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [63:0] _GEN_3661 = _T_623 ? _GEN_3633 : _GEN_3501; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire  _GEN_3663 = _T_623 ? _GEN_3635 : _GEN_3503; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [63:0] _GEN_3664 = _T_623 ? _GEN_3636 : _GEN_3504; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [63:0] _GEN_3670 = _T_623 ? _GEN_3642 : _GEN_3510; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire  _GEN_3672 = _T_623 ? _GEN_3644 : _GEN_3512; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [6:0] _GEN_3673 = _T_623 ? _GEN_3645 : _GEN_3513; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire [63:0] _GEN_3674 = _T_623 ? _GEN_3646 : _GEN_3514; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 337:20]
  wire  _GEN_3684 = _T_699 | _GEN_3672; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 346:24 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_3691 = 2'h3 == io_now_internal_privilegeMode | (2'h1 == io_now_internal_privilegeMode | (2'h0 ==
    io_now_internal_privilegeMode | _GEN_3684)); // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 354:42 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_3702 = _T_705 ? _GEN_3691 : _GEN_3684; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 352:23]
  wire  next_reg_signBit_3 = _T_844[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_346 = next_reg_signBit_3 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_347 = {_next_reg_T_346,_T_844[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_3713 = 5'h1 == rd ? _next_reg_T_347 : _GEN_3182; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3714 = 5'h2 == rd ? _next_reg_T_347 : _GEN_3183; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3715 = 5'h3 == rd ? _next_reg_T_347 : _GEN_3184; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3716 = 5'h4 == rd ? _next_reg_T_347 : _GEN_3185; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3717 = 5'h5 == rd ? _next_reg_T_347 : _GEN_3186; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3718 = 5'h6 == rd ? _next_reg_T_347 : _GEN_3187; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3719 = 5'h7 == rd ? _next_reg_T_347 : _GEN_3188; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3720 = 5'h8 == rd ? _next_reg_T_347 : _GEN_3189; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3721 = 5'h9 == rd ? _next_reg_T_347 : _GEN_3190; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3722 = 5'ha == rd ? _next_reg_T_347 : _GEN_3191; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3723 = 5'hb == rd ? _next_reg_T_347 : _GEN_3192; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3724 = 5'hc == rd ? _next_reg_T_347 : _GEN_3193; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3725 = 5'hd == rd ? _next_reg_T_347 : _GEN_3194; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3726 = 5'he == rd ? _next_reg_T_347 : _GEN_3195; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3727 = 5'hf == rd ? _next_reg_T_347 : _GEN_3196; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3728 = 5'h10 == rd ? _next_reg_T_347 : _GEN_3197; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3729 = 5'h11 == rd ? _next_reg_T_347 : _GEN_3198; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3730 = 5'h12 == rd ? _next_reg_T_347 : _GEN_3199; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3731 = 5'h13 == rd ? _next_reg_T_347 : _GEN_3200; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3732 = 5'h14 == rd ? _next_reg_T_347 : _GEN_3201; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3733 = 5'h15 == rd ? _next_reg_T_347 : _GEN_3202; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3734 = 5'h16 == rd ? _next_reg_T_347 : _GEN_3203; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3735 = 5'h17 == rd ? _next_reg_T_347 : _GEN_3204; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3736 = 5'h18 == rd ? _next_reg_T_347 : _GEN_3205; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3737 = 5'h19 == rd ? _next_reg_T_347 : _GEN_3206; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3738 = 5'h1a == rd ? _next_reg_T_347 : _GEN_3207; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3739 = 5'h1b == rd ? _next_reg_T_347 : _GEN_3208; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3740 = 5'h1c == rd ? _next_reg_T_347 : _GEN_3209; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3741 = 5'h1d == rd ? _next_reg_T_347 : _GEN_3210; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3742 = 5'h1e == rd ? _next_reg_T_347 : _GEN_3211; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3743 = 5'h1f == rd ? _next_reg_T_347 : _GEN_3212; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:{47,47}]
  wire [63:0] _GEN_3752 = _T_720 ? _GEN_3713 : _GEN_3182; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3753 = _T_720 ? _GEN_3714 : _GEN_3183; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3754 = _T_720 ? _GEN_3715 : _GEN_3184; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3755 = _T_720 ? _GEN_3716 : _GEN_3185; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3756 = _T_720 ? _GEN_3717 : _GEN_3186; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3757 = _T_720 ? _GEN_3718 : _GEN_3187; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3758 = _T_720 ? _GEN_3719 : _GEN_3188; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3759 = _T_720 ? _GEN_3720 : _GEN_3189; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3760 = _T_720 ? _GEN_3721 : _GEN_3190; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3761 = _T_720 ? _GEN_3722 : _GEN_3191; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3762 = _T_720 ? _GEN_3723 : _GEN_3192; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3763 = _T_720 ? _GEN_3724 : _GEN_3193; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3764 = _T_720 ? _GEN_3725 : _GEN_3194; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3765 = _T_720 ? _GEN_3726 : _GEN_3195; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3766 = _T_720 ? _GEN_3727 : _GEN_3196; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3767 = _T_720 ? _GEN_3728 : _GEN_3197; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3768 = _T_720 ? _GEN_3729 : _GEN_3198; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3769 = _T_720 ? _GEN_3730 : _GEN_3199; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3770 = _T_720 ? _GEN_3731 : _GEN_3200; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3771 = _T_720 ? _GEN_3732 : _GEN_3201; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3772 = _T_720 ? _GEN_3733 : _GEN_3202; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3773 = _T_720 ? _GEN_3734 : _GEN_3203; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3774 = _T_720 ? _GEN_3735 : _GEN_3204; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3775 = _T_720 ? _GEN_3736 : _GEN_3205; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3776 = _T_720 ? _GEN_3737 : _GEN_3206; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3777 = _T_720 ? _GEN_3738 : _GEN_3207; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3778 = _T_720 ? _GEN_3739 : _GEN_3208; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3779 = _T_720 ? _GEN_3740 : _GEN_3209; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3780 = _T_720 ? _GEN_3741 : _GEN_3210; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3781 = _T_720 ? _GEN_3742 : _GEN_3211; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [63:0] _GEN_3782 = _T_720 ? _GEN_3743 : _GEN_3212; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 381:23]
  wire [126:0] _GEN_2 = {{63'd0}, _GEN_101}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:62]
  wire [126:0] _next_reg_T_349 = _GEN_2 << imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:62]
  wire [63:0] _GEN_3784 = 5'h1 == rd ? _next_reg_T_349[63:0] : _GEN_3752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3785 = 5'h2 == rd ? _next_reg_T_349[63:0] : _GEN_3753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3786 = 5'h3 == rd ? _next_reg_T_349[63:0] : _GEN_3754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3787 = 5'h4 == rd ? _next_reg_T_349[63:0] : _GEN_3755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3788 = 5'h5 == rd ? _next_reg_T_349[63:0] : _GEN_3756; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3789 = 5'h6 == rd ? _next_reg_T_349[63:0] : _GEN_3757; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3790 = 5'h7 == rd ? _next_reg_T_349[63:0] : _GEN_3758; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3791 = 5'h8 == rd ? _next_reg_T_349[63:0] : _GEN_3759; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3792 = 5'h9 == rd ? _next_reg_T_349[63:0] : _GEN_3760; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3793 = 5'ha == rd ? _next_reg_T_349[63:0] : _GEN_3761; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3794 = 5'hb == rd ? _next_reg_T_349[63:0] : _GEN_3762; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3795 = 5'hc == rd ? _next_reg_T_349[63:0] : _GEN_3763; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3796 = 5'hd == rd ? _next_reg_T_349[63:0] : _GEN_3764; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3797 = 5'he == rd ? _next_reg_T_349[63:0] : _GEN_3765; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3798 = 5'hf == rd ? _next_reg_T_349[63:0] : _GEN_3766; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3799 = 5'h10 == rd ? _next_reg_T_349[63:0] : _GEN_3767; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3800 = 5'h11 == rd ? _next_reg_T_349[63:0] : _GEN_3768; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3801 = 5'h12 == rd ? _next_reg_T_349[63:0] : _GEN_3769; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3802 = 5'h13 == rd ? _next_reg_T_349[63:0] : _GEN_3770; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3803 = 5'h14 == rd ? _next_reg_T_349[63:0] : _GEN_3771; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3804 = 5'h15 == rd ? _next_reg_T_349[63:0] : _GEN_3772; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3805 = 5'h16 == rd ? _next_reg_T_349[63:0] : _GEN_3773; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3806 = 5'h17 == rd ? _next_reg_T_349[63:0] : _GEN_3774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3807 = 5'h18 == rd ? _next_reg_T_349[63:0] : _GEN_3775; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3808 = 5'h19 == rd ? _next_reg_T_349[63:0] : _GEN_3776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3809 = 5'h1a == rd ? _next_reg_T_349[63:0] : _GEN_3777; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3810 = 5'h1b == rd ? _next_reg_T_349[63:0] : _GEN_3778; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3811 = 5'h1c == rd ? _next_reg_T_349[63:0] : _GEN_3779; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3812 = 5'h1d == rd ? _next_reg_T_349[63:0] : _GEN_3780; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3813 = 5'h1e == rd ? _next_reg_T_349[63:0] : _GEN_3781; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3814 = 5'h1f == rd ? _next_reg_T_349[63:0] : _GEN_3782; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:{46,46}]
  wire [63:0] _GEN_3823 = _T_726 ? _GEN_3784 : _GEN_3752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3824 = _T_726 ? _GEN_3785 : _GEN_3753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3825 = _T_726 ? _GEN_3786 : _GEN_3754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3826 = _T_726 ? _GEN_3787 : _GEN_3755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3827 = _T_726 ? _GEN_3788 : _GEN_3756; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3828 = _T_726 ? _GEN_3789 : _GEN_3757; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3829 = _T_726 ? _GEN_3790 : _GEN_3758; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3830 = _T_726 ? _GEN_3791 : _GEN_3759; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3831 = _T_726 ? _GEN_3792 : _GEN_3760; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3832 = _T_726 ? _GEN_3793 : _GEN_3761; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3833 = _T_726 ? _GEN_3794 : _GEN_3762; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3834 = _T_726 ? _GEN_3795 : _GEN_3763; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3835 = _T_726 ? _GEN_3796 : _GEN_3764; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3836 = _T_726 ? _GEN_3797 : _GEN_3765; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3837 = _T_726 ? _GEN_3798 : _GEN_3766; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3838 = _T_726 ? _GEN_3799 : _GEN_3767; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3839 = _T_726 ? _GEN_3800 : _GEN_3768; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3840 = _T_726 ? _GEN_3801 : _GEN_3769; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3841 = _T_726 ? _GEN_3802 : _GEN_3770; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3842 = _T_726 ? _GEN_3803 : _GEN_3771; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3843 = _T_726 ? _GEN_3804 : _GEN_3772; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3844 = _T_726 ? _GEN_3805 : _GEN_3773; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3845 = _T_726 ? _GEN_3806 : _GEN_3774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3846 = _T_726 ? _GEN_3807 : _GEN_3775; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3847 = _T_726 ? _GEN_3808 : _GEN_3776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3848 = _T_726 ? _GEN_3809 : _GEN_3777; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3849 = _T_726 ? _GEN_3810 : _GEN_3778; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3850 = _T_726 ? _GEN_3811 : _GEN_3779; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3851 = _T_726 ? _GEN_3812 : _GEN_3780; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3852 = _T_726 ? _GEN_3813 : _GEN_3781; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _GEN_3853 = _T_726 ? _GEN_3814 : _GEN_3782; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 383:22]
  wire [63:0] _next_reg_T_351 = _GEN_101 >> imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:62]
  wire [63:0] _GEN_3855 = 5'h1 == rd ? _next_reg_T_351 : _GEN_3823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3856 = 5'h2 == rd ? _next_reg_T_351 : _GEN_3824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3857 = 5'h3 == rd ? _next_reg_T_351 : _GEN_3825; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3858 = 5'h4 == rd ? _next_reg_T_351 : _GEN_3826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3859 = 5'h5 == rd ? _next_reg_T_351 : _GEN_3827; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3860 = 5'h6 == rd ? _next_reg_T_351 : _GEN_3828; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3861 = 5'h7 == rd ? _next_reg_T_351 : _GEN_3829; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3862 = 5'h8 == rd ? _next_reg_T_351 : _GEN_3830; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3863 = 5'h9 == rd ? _next_reg_T_351 : _GEN_3831; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3864 = 5'ha == rd ? _next_reg_T_351 : _GEN_3832; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3865 = 5'hb == rd ? _next_reg_T_351 : _GEN_3833; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3866 = 5'hc == rd ? _next_reg_T_351 : _GEN_3834; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3867 = 5'hd == rd ? _next_reg_T_351 : _GEN_3835; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3868 = 5'he == rd ? _next_reg_T_351 : _GEN_3836; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3869 = 5'hf == rd ? _next_reg_T_351 : _GEN_3837; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3870 = 5'h10 == rd ? _next_reg_T_351 : _GEN_3838; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3871 = 5'h11 == rd ? _next_reg_T_351 : _GEN_3839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3872 = 5'h12 == rd ? _next_reg_T_351 : _GEN_3840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3873 = 5'h13 == rd ? _next_reg_T_351 : _GEN_3841; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3874 = 5'h14 == rd ? _next_reg_T_351 : _GEN_3842; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3875 = 5'h15 == rd ? _next_reg_T_351 : _GEN_3843; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3876 = 5'h16 == rd ? _next_reg_T_351 : _GEN_3844; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3877 = 5'h17 == rd ? _next_reg_T_351 : _GEN_3845; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3878 = 5'h18 == rd ? _next_reg_T_351 : _GEN_3846; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3879 = 5'h19 == rd ? _next_reg_T_351 : _GEN_3847; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3880 = 5'h1a == rd ? _next_reg_T_351 : _GEN_3848; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3881 = 5'h1b == rd ? _next_reg_T_351 : _GEN_3849; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3882 = 5'h1c == rd ? _next_reg_T_351 : _GEN_3850; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3883 = 5'h1d == rd ? _next_reg_T_351 : _GEN_3851; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3884 = 5'h1e == rd ? _next_reg_T_351 : _GEN_3852; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3885 = 5'h1f == rd ? _next_reg_T_351 : _GEN_3853; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:{46,46}]
  wire [63:0] _GEN_3894 = _T_732 ? _GEN_3855 : _GEN_3823; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3895 = _T_732 ? _GEN_3856 : _GEN_3824; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3896 = _T_732 ? _GEN_3857 : _GEN_3825; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3897 = _T_732 ? _GEN_3858 : _GEN_3826; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3898 = _T_732 ? _GEN_3859 : _GEN_3827; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3899 = _T_732 ? _GEN_3860 : _GEN_3828; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3900 = _T_732 ? _GEN_3861 : _GEN_3829; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3901 = _T_732 ? _GEN_3862 : _GEN_3830; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3902 = _T_732 ? _GEN_3863 : _GEN_3831; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3903 = _T_732 ? _GEN_3864 : _GEN_3832; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3904 = _T_732 ? _GEN_3865 : _GEN_3833; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3905 = _T_732 ? _GEN_3866 : _GEN_3834; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3906 = _T_732 ? _GEN_3867 : _GEN_3835; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3907 = _T_732 ? _GEN_3868 : _GEN_3836; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3908 = _T_732 ? _GEN_3869 : _GEN_3837; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3909 = _T_732 ? _GEN_3870 : _GEN_3838; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3910 = _T_732 ? _GEN_3871 : _GEN_3839; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3911 = _T_732 ? _GEN_3872 : _GEN_3840; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3912 = _T_732 ? _GEN_3873 : _GEN_3841; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3913 = _T_732 ? _GEN_3874 : _GEN_3842; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3914 = _T_732 ? _GEN_3875 : _GEN_3843; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3915 = _T_732 ? _GEN_3876 : _GEN_3844; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3916 = _T_732 ? _GEN_3877 : _GEN_3845; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3917 = _T_732 ? _GEN_3878 : _GEN_3846; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3918 = _T_732 ? _GEN_3879 : _GEN_3847; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3919 = _T_732 ? _GEN_3880 : _GEN_3848; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3920 = _T_732 ? _GEN_3881 : _GEN_3849; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3921 = _T_732 ? _GEN_3882 : _GEN_3850; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3922 = _T_732 ? _GEN_3883 : _GEN_3851; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3923 = _T_732 ? _GEN_3884 : _GEN_3852; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _GEN_3924 = _T_732 ? _GEN_3885 : _GEN_3853; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 384:22]
  wire [63:0] _next_reg_T_355 = $signed(_T_325) >>> imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:84]
  wire [63:0] _GEN_3926 = 5'h1 == rd ? _next_reg_T_355 : _GEN_3894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3927 = 5'h2 == rd ? _next_reg_T_355 : _GEN_3895; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3928 = 5'h3 == rd ? _next_reg_T_355 : _GEN_3896; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3929 = 5'h4 == rd ? _next_reg_T_355 : _GEN_3897; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3930 = 5'h5 == rd ? _next_reg_T_355 : _GEN_3898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3931 = 5'h6 == rd ? _next_reg_T_355 : _GEN_3899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3932 = 5'h7 == rd ? _next_reg_T_355 : _GEN_3900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3933 = 5'h8 == rd ? _next_reg_T_355 : _GEN_3901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3934 = 5'h9 == rd ? _next_reg_T_355 : _GEN_3902; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3935 = 5'ha == rd ? _next_reg_T_355 : _GEN_3903; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3936 = 5'hb == rd ? _next_reg_T_355 : _GEN_3904; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3937 = 5'hc == rd ? _next_reg_T_355 : _GEN_3905; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3938 = 5'hd == rd ? _next_reg_T_355 : _GEN_3906; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3939 = 5'he == rd ? _next_reg_T_355 : _GEN_3907; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3940 = 5'hf == rd ? _next_reg_T_355 : _GEN_3908; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3941 = 5'h10 == rd ? _next_reg_T_355 : _GEN_3909; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3942 = 5'h11 == rd ? _next_reg_T_355 : _GEN_3910; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3943 = 5'h12 == rd ? _next_reg_T_355 : _GEN_3911; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3944 = 5'h13 == rd ? _next_reg_T_355 : _GEN_3912; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3945 = 5'h14 == rd ? _next_reg_T_355 : _GEN_3913; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3946 = 5'h15 == rd ? _next_reg_T_355 : _GEN_3914; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3947 = 5'h16 == rd ? _next_reg_T_355 : _GEN_3915; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3948 = 5'h17 == rd ? _next_reg_T_355 : _GEN_3916; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3949 = 5'h18 == rd ? _next_reg_T_355 : _GEN_3917; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3950 = 5'h19 == rd ? _next_reg_T_355 : _GEN_3918; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3951 = 5'h1a == rd ? _next_reg_T_355 : _GEN_3919; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3952 = 5'h1b == rd ? _next_reg_T_355 : _GEN_3920; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3953 = 5'h1c == rd ? _next_reg_T_355 : _GEN_3921; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3954 = 5'h1d == rd ? _next_reg_T_355 : _GEN_3922; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3955 = 5'h1e == rd ? _next_reg_T_355 : _GEN_3923; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3956 = 5'h1f == rd ? _next_reg_T_355 : _GEN_3924; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:{46,46}]
  wire [63:0] _GEN_3965 = _T_738 ? _GEN_3926 : _GEN_3894; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3966 = _T_738 ? _GEN_3927 : _GEN_3895; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3967 = _T_738 ? _GEN_3928 : _GEN_3896; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3968 = _T_738 ? _GEN_3929 : _GEN_3897; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3969 = _T_738 ? _GEN_3930 : _GEN_3898; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3970 = _T_738 ? _GEN_3931 : _GEN_3899; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3971 = _T_738 ? _GEN_3932 : _GEN_3900; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3972 = _T_738 ? _GEN_3933 : _GEN_3901; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3973 = _T_738 ? _GEN_3934 : _GEN_3902; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3974 = _T_738 ? _GEN_3935 : _GEN_3903; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3975 = _T_738 ? _GEN_3936 : _GEN_3904; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3976 = _T_738 ? _GEN_3937 : _GEN_3905; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3977 = _T_738 ? _GEN_3938 : _GEN_3906; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3978 = _T_738 ? _GEN_3939 : _GEN_3907; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3979 = _T_738 ? _GEN_3940 : _GEN_3908; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3980 = _T_738 ? _GEN_3941 : _GEN_3909; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3981 = _T_738 ? _GEN_3942 : _GEN_3910; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3982 = _T_738 ? _GEN_3943 : _GEN_3911; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3983 = _T_738 ? _GEN_3944 : _GEN_3912; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3984 = _T_738 ? _GEN_3945 : _GEN_3913; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3985 = _T_738 ? _GEN_3946 : _GEN_3914; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3986 = _T_738 ? _GEN_3947 : _GEN_3915; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3987 = _T_738 ? _GEN_3948 : _GEN_3916; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3988 = _T_738 ? _GEN_3949 : _GEN_3917; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3989 = _T_738 ? _GEN_3950 : _GEN_3918; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3990 = _T_738 ? _GEN_3951 : _GEN_3919; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3991 = _T_738 ? _GEN_3952 : _GEN_3920; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3992 = _T_738 ? _GEN_3953 : _GEN_3921; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3993 = _T_738 ? _GEN_3954 : _GEN_3922; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3994 = _T_738 ? _GEN_3955 : _GEN_3923; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [63:0] _GEN_3995 = _T_738 ? _GEN_3956 : _GEN_3924; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 385:22]
  wire [62:0] _GEN_3 = {{31'd0}, _GEN_101[31:0]}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:79]
  wire [62:0] _next_reg_T_358 = _GEN_3 << imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:79]
  wire  next_reg_signBit_4 = _next_reg_T_358[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_361 = next_reg_signBit_4 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_362 = {_next_reg_T_361,_next_reg_T_358[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_3997 = 5'h1 == rd ? _next_reg_T_362 : _GEN_3965; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_3998 = 5'h2 == rd ? _next_reg_T_362 : _GEN_3966; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_3999 = 5'h3 == rd ? _next_reg_T_362 : _GEN_3967; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4000 = 5'h4 == rd ? _next_reg_T_362 : _GEN_3968; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4001 = 5'h5 == rd ? _next_reg_T_362 : _GEN_3969; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4002 = 5'h6 == rd ? _next_reg_T_362 : _GEN_3970; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4003 = 5'h7 == rd ? _next_reg_T_362 : _GEN_3971; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4004 = 5'h8 == rd ? _next_reg_T_362 : _GEN_3972; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4005 = 5'h9 == rd ? _next_reg_T_362 : _GEN_3973; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4006 = 5'ha == rd ? _next_reg_T_362 : _GEN_3974; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4007 = 5'hb == rd ? _next_reg_T_362 : _GEN_3975; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4008 = 5'hc == rd ? _next_reg_T_362 : _GEN_3976; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4009 = 5'hd == rd ? _next_reg_T_362 : _GEN_3977; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4010 = 5'he == rd ? _next_reg_T_362 : _GEN_3978; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4011 = 5'hf == rd ? _next_reg_T_362 : _GEN_3979; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4012 = 5'h10 == rd ? _next_reg_T_362 : _GEN_3980; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4013 = 5'h11 == rd ? _next_reg_T_362 : _GEN_3981; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4014 = 5'h12 == rd ? _next_reg_T_362 : _GEN_3982; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4015 = 5'h13 == rd ? _next_reg_T_362 : _GEN_3983; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4016 = 5'h14 == rd ? _next_reg_T_362 : _GEN_3984; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4017 = 5'h15 == rd ? _next_reg_T_362 : _GEN_3985; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4018 = 5'h16 == rd ? _next_reg_T_362 : _GEN_3986; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4019 = 5'h17 == rd ? _next_reg_T_362 : _GEN_3987; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4020 = 5'h18 == rd ? _next_reg_T_362 : _GEN_3988; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4021 = 5'h19 == rd ? _next_reg_T_362 : _GEN_3989; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4022 = 5'h1a == rd ? _next_reg_T_362 : _GEN_3990; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4023 = 5'h1b == rd ? _next_reg_T_362 : _GEN_3991; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4024 = 5'h1c == rd ? _next_reg_T_362 : _GEN_3992; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4025 = 5'h1d == rd ? _next_reg_T_362 : _GEN_3993; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4026 = 5'h1e == rd ? _next_reg_T_362 : _GEN_3994; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4027 = 5'h1f == rd ? _next_reg_T_362 : _GEN_3995; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:{47,47}]
  wire [63:0] _GEN_4036 = _T_744 ? _GEN_3997 : _GEN_3965; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4037 = _T_744 ? _GEN_3998 : _GEN_3966; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4038 = _T_744 ? _GEN_3999 : _GEN_3967; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4039 = _T_744 ? _GEN_4000 : _GEN_3968; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4040 = _T_744 ? _GEN_4001 : _GEN_3969; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4041 = _T_744 ? _GEN_4002 : _GEN_3970; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4042 = _T_744 ? _GEN_4003 : _GEN_3971; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4043 = _T_744 ? _GEN_4004 : _GEN_3972; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4044 = _T_744 ? _GEN_4005 : _GEN_3973; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4045 = _T_744 ? _GEN_4006 : _GEN_3974; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4046 = _T_744 ? _GEN_4007 : _GEN_3975; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4047 = _T_744 ? _GEN_4008 : _GEN_3976; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4048 = _T_744 ? _GEN_4009 : _GEN_3977; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4049 = _T_744 ? _GEN_4010 : _GEN_3978; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4050 = _T_744 ? _GEN_4011 : _GEN_3979; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4051 = _T_744 ? _GEN_4012 : _GEN_3980; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4052 = _T_744 ? _GEN_4013 : _GEN_3981; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4053 = _T_744 ? _GEN_4014 : _GEN_3982; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4054 = _T_744 ? _GEN_4015 : _GEN_3983; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4055 = _T_744 ? _GEN_4016 : _GEN_3984; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4056 = _T_744 ? _GEN_4017 : _GEN_3985; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4057 = _T_744 ? _GEN_4018 : _GEN_3986; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4058 = _T_744 ? _GEN_4019 : _GEN_3987; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4059 = _T_744 ? _GEN_4020 : _GEN_3988; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4060 = _T_744 ? _GEN_4021 : _GEN_3989; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4061 = _T_744 ? _GEN_4022 : _GEN_3990; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4062 = _T_744 ? _GEN_4023 : _GEN_3991; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4063 = _T_744 ? _GEN_4024 : _GEN_3992; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4064 = _T_744 ? _GEN_4025 : _GEN_3993; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4065 = _T_744 ? _GEN_4026 : _GEN_3994; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [63:0] _GEN_4066 = _T_744 ? _GEN_4027 : _GEN_3995; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 387:23]
  wire [31:0] _next_reg_T_365 = _GEN_101[31:0] >> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:78]
  wire  next_reg_signBit_5 = _next_reg_T_365[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_367 = next_reg_signBit_5 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_368 = {_next_reg_T_367,_next_reg_T_365}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_4068 = 5'h1 == rd ? _next_reg_T_368 : _GEN_4036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4069 = 5'h2 == rd ? _next_reg_T_368 : _GEN_4037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4070 = 5'h3 == rd ? _next_reg_T_368 : _GEN_4038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4071 = 5'h4 == rd ? _next_reg_T_368 : _GEN_4039; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4072 = 5'h5 == rd ? _next_reg_T_368 : _GEN_4040; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4073 = 5'h6 == rd ? _next_reg_T_368 : _GEN_4041; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4074 = 5'h7 == rd ? _next_reg_T_368 : _GEN_4042; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4075 = 5'h8 == rd ? _next_reg_T_368 : _GEN_4043; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4076 = 5'h9 == rd ? _next_reg_T_368 : _GEN_4044; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4077 = 5'ha == rd ? _next_reg_T_368 : _GEN_4045; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4078 = 5'hb == rd ? _next_reg_T_368 : _GEN_4046; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4079 = 5'hc == rd ? _next_reg_T_368 : _GEN_4047; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4080 = 5'hd == rd ? _next_reg_T_368 : _GEN_4048; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4081 = 5'he == rd ? _next_reg_T_368 : _GEN_4049; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4082 = 5'hf == rd ? _next_reg_T_368 : _GEN_4050; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4083 = 5'h10 == rd ? _next_reg_T_368 : _GEN_4051; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4084 = 5'h11 == rd ? _next_reg_T_368 : _GEN_4052; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4085 = 5'h12 == rd ? _next_reg_T_368 : _GEN_4053; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4086 = 5'h13 == rd ? _next_reg_T_368 : _GEN_4054; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4087 = 5'h14 == rd ? _next_reg_T_368 : _GEN_4055; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4088 = 5'h15 == rd ? _next_reg_T_368 : _GEN_4056; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4089 = 5'h16 == rd ? _next_reg_T_368 : _GEN_4057; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4090 = 5'h17 == rd ? _next_reg_T_368 : _GEN_4058; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4091 = 5'h18 == rd ? _next_reg_T_368 : _GEN_4059; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4092 = 5'h19 == rd ? _next_reg_T_368 : _GEN_4060; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4093 = 5'h1a == rd ? _next_reg_T_368 : _GEN_4061; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4094 = 5'h1b == rd ? _next_reg_T_368 : _GEN_4062; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4095 = 5'h1c == rd ? _next_reg_T_368 : _GEN_4063; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4096 = 5'h1d == rd ? _next_reg_T_368 : _GEN_4064; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4097 = 5'h1e == rd ? _next_reg_T_368 : _GEN_4065; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4098 = 5'h1f == rd ? _next_reg_T_368 : _GEN_4066; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:{47,47}]
  wire [63:0] _GEN_4107 = _T_750 ? _GEN_4068 : _GEN_4036; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4108 = _T_750 ? _GEN_4069 : _GEN_4037; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4109 = _T_750 ? _GEN_4070 : _GEN_4038; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4110 = _T_750 ? _GEN_4071 : _GEN_4039; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4111 = _T_750 ? _GEN_4072 : _GEN_4040; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4112 = _T_750 ? _GEN_4073 : _GEN_4041; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4113 = _T_750 ? _GEN_4074 : _GEN_4042; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4114 = _T_750 ? _GEN_4075 : _GEN_4043; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4115 = _T_750 ? _GEN_4076 : _GEN_4044; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4116 = _T_750 ? _GEN_4077 : _GEN_4045; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4117 = _T_750 ? _GEN_4078 : _GEN_4046; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4118 = _T_750 ? _GEN_4079 : _GEN_4047; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4119 = _T_750 ? _GEN_4080 : _GEN_4048; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4120 = _T_750 ? _GEN_4081 : _GEN_4049; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4121 = _T_750 ? _GEN_4082 : _GEN_4050; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4122 = _T_750 ? _GEN_4083 : _GEN_4051; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4123 = _T_750 ? _GEN_4084 : _GEN_4052; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4124 = _T_750 ? _GEN_4085 : _GEN_4053; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4125 = _T_750 ? _GEN_4086 : _GEN_4054; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4126 = _T_750 ? _GEN_4087 : _GEN_4055; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4127 = _T_750 ? _GEN_4088 : _GEN_4056; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4128 = _T_750 ? _GEN_4089 : _GEN_4057; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4129 = _T_750 ? _GEN_4090 : _GEN_4058; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4130 = _T_750 ? _GEN_4091 : _GEN_4059; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4131 = _T_750 ? _GEN_4092 : _GEN_4060; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4132 = _T_750 ? _GEN_4093 : _GEN_4061; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4133 = _T_750 ? _GEN_4094 : _GEN_4062; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4134 = _T_750 ? _GEN_4095 : _GEN_4063; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4135 = _T_750 ? _GEN_4096 : _GEN_4064; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4136 = _T_750 ? _GEN_4097 : _GEN_4065; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [63:0] _GEN_4137 = _T_750 ? _GEN_4098 : _GEN_4066; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 388:23]
  wire [31:0] _next_reg_T_370 = _GEN_101[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:79]
  wire [31:0] _next_reg_T_373 = $signed(_next_reg_T_370) >>> imm[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:100]
  wire  next_reg_signBit_6 = _next_reg_T_373[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_375 = next_reg_signBit_6 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_376 = {_next_reg_T_375,_next_reg_T_373}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_4139 = 5'h1 == rd ? _next_reg_T_376 : _GEN_4107; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4140 = 5'h2 == rd ? _next_reg_T_376 : _GEN_4108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4141 = 5'h3 == rd ? _next_reg_T_376 : _GEN_4109; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4142 = 5'h4 == rd ? _next_reg_T_376 : _GEN_4110; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4143 = 5'h5 == rd ? _next_reg_T_376 : _GEN_4111; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4144 = 5'h6 == rd ? _next_reg_T_376 : _GEN_4112; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4145 = 5'h7 == rd ? _next_reg_T_376 : _GEN_4113; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4146 = 5'h8 == rd ? _next_reg_T_376 : _GEN_4114; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4147 = 5'h9 == rd ? _next_reg_T_376 : _GEN_4115; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4148 = 5'ha == rd ? _next_reg_T_376 : _GEN_4116; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4149 = 5'hb == rd ? _next_reg_T_376 : _GEN_4117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4150 = 5'hc == rd ? _next_reg_T_376 : _GEN_4118; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4151 = 5'hd == rd ? _next_reg_T_376 : _GEN_4119; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4152 = 5'he == rd ? _next_reg_T_376 : _GEN_4120; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4153 = 5'hf == rd ? _next_reg_T_376 : _GEN_4121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4154 = 5'h10 == rd ? _next_reg_T_376 : _GEN_4122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4155 = 5'h11 == rd ? _next_reg_T_376 : _GEN_4123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4156 = 5'h12 == rd ? _next_reg_T_376 : _GEN_4124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4157 = 5'h13 == rd ? _next_reg_T_376 : _GEN_4125; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4158 = 5'h14 == rd ? _next_reg_T_376 : _GEN_4126; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4159 = 5'h15 == rd ? _next_reg_T_376 : _GEN_4127; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4160 = 5'h16 == rd ? _next_reg_T_376 : _GEN_4128; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4161 = 5'h17 == rd ? _next_reg_T_376 : _GEN_4129; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4162 = 5'h18 == rd ? _next_reg_T_376 : _GEN_4130; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4163 = 5'h19 == rd ? _next_reg_T_376 : _GEN_4131; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4164 = 5'h1a == rd ? _next_reg_T_376 : _GEN_4132; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4165 = 5'h1b == rd ? _next_reg_T_376 : _GEN_4133; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4166 = 5'h1c == rd ? _next_reg_T_376 : _GEN_4134; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4167 = 5'h1d == rd ? _next_reg_T_376 : _GEN_4135; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4168 = 5'h1e == rd ? _next_reg_T_376 : _GEN_4136; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4169 = 5'h1f == rd ? _next_reg_T_376 : _GEN_4137; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:{47,47}]
  wire [63:0] _GEN_4178 = _T_756 ? _GEN_4139 : _GEN_4107; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4179 = _T_756 ? _GEN_4140 : _GEN_4108; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4180 = _T_756 ? _GEN_4141 : _GEN_4109; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4181 = _T_756 ? _GEN_4142 : _GEN_4110; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4182 = _T_756 ? _GEN_4143 : _GEN_4111; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4183 = _T_756 ? _GEN_4144 : _GEN_4112; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4184 = _T_756 ? _GEN_4145 : _GEN_4113; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4185 = _T_756 ? _GEN_4146 : _GEN_4114; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4186 = _T_756 ? _GEN_4147 : _GEN_4115; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4187 = _T_756 ? _GEN_4148 : _GEN_4116; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4188 = _T_756 ? _GEN_4149 : _GEN_4117; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4189 = _T_756 ? _GEN_4150 : _GEN_4118; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4190 = _T_756 ? _GEN_4151 : _GEN_4119; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4191 = _T_756 ? _GEN_4152 : _GEN_4120; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4192 = _T_756 ? _GEN_4153 : _GEN_4121; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4193 = _T_756 ? _GEN_4154 : _GEN_4122; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4194 = _T_756 ? _GEN_4155 : _GEN_4123; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4195 = _T_756 ? _GEN_4156 : _GEN_4124; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4196 = _T_756 ? _GEN_4157 : _GEN_4125; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4197 = _T_756 ? _GEN_4158 : _GEN_4126; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4198 = _T_756 ? _GEN_4159 : _GEN_4127; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4199 = _T_756 ? _GEN_4160 : _GEN_4128; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4200 = _T_756 ? _GEN_4161 : _GEN_4129; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4201 = _T_756 ? _GEN_4162 : _GEN_4130; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4202 = _T_756 ? _GEN_4163 : _GEN_4131; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4203 = _T_756 ? _GEN_4164 : _GEN_4132; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4204 = _T_756 ? _GEN_4165 : _GEN_4133; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4205 = _T_756 ? _GEN_4166 : _GEN_4134; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4206 = _T_756 ? _GEN_4167 : _GEN_4135; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4207 = _T_756 ? _GEN_4168 : _GEN_4136; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [63:0] _GEN_4208 = _T_756 ? _GEN_4169 : _GEN_4137; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 389:23]
  wire [126:0] _GEN_4 = {{63'd0}, _GEN_101}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:61]
  wire [126:0] _next_reg_T_378 = _GEN_4 << _GEN_910[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:61]
  wire [63:0] _GEN_4210 = 5'h1 == rd ? _next_reg_T_378[63:0] : _GEN_4178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4211 = 5'h2 == rd ? _next_reg_T_378[63:0] : _GEN_4179; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4212 = 5'h3 == rd ? _next_reg_T_378[63:0] : _GEN_4180; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4213 = 5'h4 == rd ? _next_reg_T_378[63:0] : _GEN_4181; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4214 = 5'h5 == rd ? _next_reg_T_378[63:0] : _GEN_4182; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4215 = 5'h6 == rd ? _next_reg_T_378[63:0] : _GEN_4183; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4216 = 5'h7 == rd ? _next_reg_T_378[63:0] : _GEN_4184; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4217 = 5'h8 == rd ? _next_reg_T_378[63:0] : _GEN_4185; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4218 = 5'h9 == rd ? _next_reg_T_378[63:0] : _GEN_4186; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4219 = 5'ha == rd ? _next_reg_T_378[63:0] : _GEN_4187; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4220 = 5'hb == rd ? _next_reg_T_378[63:0] : _GEN_4188; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4221 = 5'hc == rd ? _next_reg_T_378[63:0] : _GEN_4189; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4222 = 5'hd == rd ? _next_reg_T_378[63:0] : _GEN_4190; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4223 = 5'he == rd ? _next_reg_T_378[63:0] : _GEN_4191; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4224 = 5'hf == rd ? _next_reg_T_378[63:0] : _GEN_4192; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4225 = 5'h10 == rd ? _next_reg_T_378[63:0] : _GEN_4193; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4226 = 5'h11 == rd ? _next_reg_T_378[63:0] : _GEN_4194; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4227 = 5'h12 == rd ? _next_reg_T_378[63:0] : _GEN_4195; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4228 = 5'h13 == rd ? _next_reg_T_378[63:0] : _GEN_4196; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4229 = 5'h14 == rd ? _next_reg_T_378[63:0] : _GEN_4197; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4230 = 5'h15 == rd ? _next_reg_T_378[63:0] : _GEN_4198; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4231 = 5'h16 == rd ? _next_reg_T_378[63:0] : _GEN_4199; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4232 = 5'h17 == rd ? _next_reg_T_378[63:0] : _GEN_4200; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4233 = 5'h18 == rd ? _next_reg_T_378[63:0] : _GEN_4201; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4234 = 5'h19 == rd ? _next_reg_T_378[63:0] : _GEN_4202; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4235 = 5'h1a == rd ? _next_reg_T_378[63:0] : _GEN_4203; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4236 = 5'h1b == rd ? _next_reg_T_378[63:0] : _GEN_4204; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4237 = 5'h1c == rd ? _next_reg_T_378[63:0] : _GEN_4205; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4238 = 5'h1d == rd ? _next_reg_T_378[63:0] : _GEN_4206; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4239 = 5'h1e == rd ? _next_reg_T_378[63:0] : _GEN_4207; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4240 = 5'h1f == rd ? _next_reg_T_378[63:0] : _GEN_4208; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:{45,45}]
  wire [63:0] _GEN_4249 = _T_762 ? _GEN_4210 : _GEN_4178; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4250 = _T_762 ? _GEN_4211 : _GEN_4179; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4251 = _T_762 ? _GEN_4212 : _GEN_4180; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4252 = _T_762 ? _GEN_4213 : _GEN_4181; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4253 = _T_762 ? _GEN_4214 : _GEN_4182; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4254 = _T_762 ? _GEN_4215 : _GEN_4183; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4255 = _T_762 ? _GEN_4216 : _GEN_4184; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4256 = _T_762 ? _GEN_4217 : _GEN_4185; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4257 = _T_762 ? _GEN_4218 : _GEN_4186; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4258 = _T_762 ? _GEN_4219 : _GEN_4187; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4259 = _T_762 ? _GEN_4220 : _GEN_4188; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4260 = _T_762 ? _GEN_4221 : _GEN_4189; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4261 = _T_762 ? _GEN_4222 : _GEN_4190; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4262 = _T_762 ? _GEN_4223 : _GEN_4191; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4263 = _T_762 ? _GEN_4224 : _GEN_4192; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4264 = _T_762 ? _GEN_4225 : _GEN_4193; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4265 = _T_762 ? _GEN_4226 : _GEN_4194; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4266 = _T_762 ? _GEN_4227 : _GEN_4195; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4267 = _T_762 ? _GEN_4228 : _GEN_4196; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4268 = _T_762 ? _GEN_4229 : _GEN_4197; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4269 = _T_762 ? _GEN_4230 : _GEN_4198; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4270 = _T_762 ? _GEN_4231 : _GEN_4199; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4271 = _T_762 ? _GEN_4232 : _GEN_4200; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4272 = _T_762 ? _GEN_4233 : _GEN_4201; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4273 = _T_762 ? _GEN_4234 : _GEN_4202; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4274 = _T_762 ? _GEN_4235 : _GEN_4203; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4275 = _T_762 ? _GEN_4236 : _GEN_4204; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4276 = _T_762 ? _GEN_4237 : _GEN_4205; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4277 = _T_762 ? _GEN_4238 : _GEN_4206; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4278 = _T_762 ? _GEN_4239 : _GEN_4207; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _GEN_4279 = _T_762 ? _GEN_4240 : _GEN_4208; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 393:21]
  wire [63:0] _next_reg_T_380 = _GEN_101 >> _GEN_910[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:61]
  wire [63:0] _GEN_4281 = 5'h1 == rd ? _next_reg_T_380 : _GEN_4249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4282 = 5'h2 == rd ? _next_reg_T_380 : _GEN_4250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4283 = 5'h3 == rd ? _next_reg_T_380 : _GEN_4251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4284 = 5'h4 == rd ? _next_reg_T_380 : _GEN_4252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4285 = 5'h5 == rd ? _next_reg_T_380 : _GEN_4253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4286 = 5'h6 == rd ? _next_reg_T_380 : _GEN_4254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4287 = 5'h7 == rd ? _next_reg_T_380 : _GEN_4255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4288 = 5'h8 == rd ? _next_reg_T_380 : _GEN_4256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4289 = 5'h9 == rd ? _next_reg_T_380 : _GEN_4257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4290 = 5'ha == rd ? _next_reg_T_380 : _GEN_4258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4291 = 5'hb == rd ? _next_reg_T_380 : _GEN_4259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4292 = 5'hc == rd ? _next_reg_T_380 : _GEN_4260; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4293 = 5'hd == rd ? _next_reg_T_380 : _GEN_4261; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4294 = 5'he == rd ? _next_reg_T_380 : _GEN_4262; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4295 = 5'hf == rd ? _next_reg_T_380 : _GEN_4263; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4296 = 5'h10 == rd ? _next_reg_T_380 : _GEN_4264; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4297 = 5'h11 == rd ? _next_reg_T_380 : _GEN_4265; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4298 = 5'h12 == rd ? _next_reg_T_380 : _GEN_4266; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4299 = 5'h13 == rd ? _next_reg_T_380 : _GEN_4267; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4300 = 5'h14 == rd ? _next_reg_T_380 : _GEN_4268; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4301 = 5'h15 == rd ? _next_reg_T_380 : _GEN_4269; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4302 = 5'h16 == rd ? _next_reg_T_380 : _GEN_4270; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4303 = 5'h17 == rd ? _next_reg_T_380 : _GEN_4271; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4304 = 5'h18 == rd ? _next_reg_T_380 : _GEN_4272; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4305 = 5'h19 == rd ? _next_reg_T_380 : _GEN_4273; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4306 = 5'h1a == rd ? _next_reg_T_380 : _GEN_4274; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4307 = 5'h1b == rd ? _next_reg_T_380 : _GEN_4275; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4308 = 5'h1c == rd ? _next_reg_T_380 : _GEN_4276; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4309 = 5'h1d == rd ? _next_reg_T_380 : _GEN_4277; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4310 = 5'h1e == rd ? _next_reg_T_380 : _GEN_4278; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4311 = 5'h1f == rd ? _next_reg_T_380 : _GEN_4279; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:{45,45}]
  wire [63:0] _GEN_4320 = _T_769 ? _GEN_4281 : _GEN_4249; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4321 = _T_769 ? _GEN_4282 : _GEN_4250; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4322 = _T_769 ? _GEN_4283 : _GEN_4251; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4323 = _T_769 ? _GEN_4284 : _GEN_4252; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4324 = _T_769 ? _GEN_4285 : _GEN_4253; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4325 = _T_769 ? _GEN_4286 : _GEN_4254; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4326 = _T_769 ? _GEN_4287 : _GEN_4255; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4327 = _T_769 ? _GEN_4288 : _GEN_4256; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4328 = _T_769 ? _GEN_4289 : _GEN_4257; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4329 = _T_769 ? _GEN_4290 : _GEN_4258; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4330 = _T_769 ? _GEN_4291 : _GEN_4259; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4331 = _T_769 ? _GEN_4292 : _GEN_4260; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4332 = _T_769 ? _GEN_4293 : _GEN_4261; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4333 = _T_769 ? _GEN_4294 : _GEN_4262; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4334 = _T_769 ? _GEN_4295 : _GEN_4263; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4335 = _T_769 ? _GEN_4296 : _GEN_4264; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4336 = _T_769 ? _GEN_4297 : _GEN_4265; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4337 = _T_769 ? _GEN_4298 : _GEN_4266; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4338 = _T_769 ? _GEN_4299 : _GEN_4267; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4339 = _T_769 ? _GEN_4300 : _GEN_4268; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4340 = _T_769 ? _GEN_4301 : _GEN_4269; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4341 = _T_769 ? _GEN_4302 : _GEN_4270; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4342 = _T_769 ? _GEN_4303 : _GEN_4271; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4343 = _T_769 ? _GEN_4304 : _GEN_4272; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4344 = _T_769 ? _GEN_4305 : _GEN_4273; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4345 = _T_769 ? _GEN_4306 : _GEN_4274; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4346 = _T_769 ? _GEN_4307 : _GEN_4275; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4347 = _T_769 ? _GEN_4308 : _GEN_4276; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4348 = _T_769 ? _GEN_4309 : _GEN_4277; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4349 = _T_769 ? _GEN_4310 : _GEN_4278; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _GEN_4350 = _T_769 ? _GEN_4311 : _GEN_4279; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 394:21]
  wire [63:0] _next_reg_T_384 = $signed(_T_325) >>> _GEN_910[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:92]
  wire [63:0] _GEN_4352 = 5'h1 == rd ? _next_reg_T_384 : _GEN_4320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4353 = 5'h2 == rd ? _next_reg_T_384 : _GEN_4321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4354 = 5'h3 == rd ? _next_reg_T_384 : _GEN_4322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4355 = 5'h4 == rd ? _next_reg_T_384 : _GEN_4323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4356 = 5'h5 == rd ? _next_reg_T_384 : _GEN_4324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4357 = 5'h6 == rd ? _next_reg_T_384 : _GEN_4325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4358 = 5'h7 == rd ? _next_reg_T_384 : _GEN_4326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4359 = 5'h8 == rd ? _next_reg_T_384 : _GEN_4327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4360 = 5'h9 == rd ? _next_reg_T_384 : _GEN_4328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4361 = 5'ha == rd ? _next_reg_T_384 : _GEN_4329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4362 = 5'hb == rd ? _next_reg_T_384 : _GEN_4330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4363 = 5'hc == rd ? _next_reg_T_384 : _GEN_4331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4364 = 5'hd == rd ? _next_reg_T_384 : _GEN_4332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4365 = 5'he == rd ? _next_reg_T_384 : _GEN_4333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4366 = 5'hf == rd ? _next_reg_T_384 : _GEN_4334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4367 = 5'h10 == rd ? _next_reg_T_384 : _GEN_4335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4368 = 5'h11 == rd ? _next_reg_T_384 : _GEN_4336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4369 = 5'h12 == rd ? _next_reg_T_384 : _GEN_4337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4370 = 5'h13 == rd ? _next_reg_T_384 : _GEN_4338; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4371 = 5'h14 == rd ? _next_reg_T_384 : _GEN_4339; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4372 = 5'h15 == rd ? _next_reg_T_384 : _GEN_4340; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4373 = 5'h16 == rd ? _next_reg_T_384 : _GEN_4341; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4374 = 5'h17 == rd ? _next_reg_T_384 : _GEN_4342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4375 = 5'h18 == rd ? _next_reg_T_384 : _GEN_4343; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4376 = 5'h19 == rd ? _next_reg_T_384 : _GEN_4344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4377 = 5'h1a == rd ? _next_reg_T_384 : _GEN_4345; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4378 = 5'h1b == rd ? _next_reg_T_384 : _GEN_4346; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4379 = 5'h1c == rd ? _next_reg_T_384 : _GEN_4347; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4380 = 5'h1d == rd ? _next_reg_T_384 : _GEN_4348; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4381 = 5'h1e == rd ? _next_reg_T_384 : _GEN_4349; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4382 = 5'h1f == rd ? _next_reg_T_384 : _GEN_4350; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:{45,45}]
  wire [63:0] _GEN_4391 = _T_776 ? _GEN_4352 : _GEN_4320; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4392 = _T_776 ? _GEN_4353 : _GEN_4321; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4393 = _T_776 ? _GEN_4354 : _GEN_4322; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4394 = _T_776 ? _GEN_4355 : _GEN_4323; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4395 = _T_776 ? _GEN_4356 : _GEN_4324; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4396 = _T_776 ? _GEN_4357 : _GEN_4325; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4397 = _T_776 ? _GEN_4358 : _GEN_4326; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4398 = _T_776 ? _GEN_4359 : _GEN_4327; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4399 = _T_776 ? _GEN_4360 : _GEN_4328; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4400 = _T_776 ? _GEN_4361 : _GEN_4329; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4401 = _T_776 ? _GEN_4362 : _GEN_4330; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4402 = _T_776 ? _GEN_4363 : _GEN_4331; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4403 = _T_776 ? _GEN_4364 : _GEN_4332; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4404 = _T_776 ? _GEN_4365 : _GEN_4333; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4405 = _T_776 ? _GEN_4366 : _GEN_4334; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4406 = _T_776 ? _GEN_4367 : _GEN_4335; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4407 = _T_776 ? _GEN_4368 : _GEN_4336; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4408 = _T_776 ? _GEN_4369 : _GEN_4337; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4409 = _T_776 ? _GEN_4370 : _GEN_4338; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4410 = _T_776 ? _GEN_4371 : _GEN_4339; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4411 = _T_776 ? _GEN_4372 : _GEN_4340; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4412 = _T_776 ? _GEN_4373 : _GEN_4341; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4413 = _T_776 ? _GEN_4374 : _GEN_4342; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4414 = _T_776 ? _GEN_4375 : _GEN_4343; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4415 = _T_776 ? _GEN_4376 : _GEN_4344; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4416 = _T_776 ? _GEN_4377 : _GEN_4345; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4417 = _T_776 ? _GEN_4378 : _GEN_4346; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4418 = _T_776 ? _GEN_4379 : _GEN_4347; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4419 = _T_776 ? _GEN_4380 : _GEN_4348; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4420 = _T_776 ? _GEN_4381 : _GEN_4349; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [63:0] _GEN_4421 = _T_776 ? _GEN_4382 : _GEN_4350; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 396:21]
  wire [31:0] _next_reg_T_388 = _GEN_101[31:0] + _GEN_910[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:78]
  wire  next_reg_signBit_7 = _next_reg_T_388[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_391 = next_reg_signBit_7 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_392 = {_next_reg_T_391,_next_reg_T_388}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_4423 = 5'h1 == rd ? _next_reg_T_392 : _GEN_4391; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4424 = 5'h2 == rd ? _next_reg_T_392 : _GEN_4392; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4425 = 5'h3 == rd ? _next_reg_T_392 : _GEN_4393; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4426 = 5'h4 == rd ? _next_reg_T_392 : _GEN_4394; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4427 = 5'h5 == rd ? _next_reg_T_392 : _GEN_4395; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4428 = 5'h6 == rd ? _next_reg_T_392 : _GEN_4396; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4429 = 5'h7 == rd ? _next_reg_T_392 : _GEN_4397; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4430 = 5'h8 == rd ? _next_reg_T_392 : _GEN_4398; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4431 = 5'h9 == rd ? _next_reg_T_392 : _GEN_4399; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4432 = 5'ha == rd ? _next_reg_T_392 : _GEN_4400; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4433 = 5'hb == rd ? _next_reg_T_392 : _GEN_4401; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4434 = 5'hc == rd ? _next_reg_T_392 : _GEN_4402; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4435 = 5'hd == rd ? _next_reg_T_392 : _GEN_4403; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4436 = 5'he == rd ? _next_reg_T_392 : _GEN_4404; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4437 = 5'hf == rd ? _next_reg_T_392 : _GEN_4405; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4438 = 5'h10 == rd ? _next_reg_T_392 : _GEN_4406; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4439 = 5'h11 == rd ? _next_reg_T_392 : _GEN_4407; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4440 = 5'h12 == rd ? _next_reg_T_392 : _GEN_4408; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4441 = 5'h13 == rd ? _next_reg_T_392 : _GEN_4409; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4442 = 5'h14 == rd ? _next_reg_T_392 : _GEN_4410; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4443 = 5'h15 == rd ? _next_reg_T_392 : _GEN_4411; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4444 = 5'h16 == rd ? _next_reg_T_392 : _GEN_4412; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4445 = 5'h17 == rd ? _next_reg_T_392 : _GEN_4413; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4446 = 5'h18 == rd ? _next_reg_T_392 : _GEN_4414; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4447 = 5'h19 == rd ? _next_reg_T_392 : _GEN_4415; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4448 = 5'h1a == rd ? _next_reg_T_392 : _GEN_4416; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4449 = 5'h1b == rd ? _next_reg_T_392 : _GEN_4417; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4450 = 5'h1c == rd ? _next_reg_T_392 : _GEN_4418; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4451 = 5'h1d == rd ? _next_reg_T_392 : _GEN_4419; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4452 = 5'h1e == rd ? _next_reg_T_392 : _GEN_4420; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4453 = 5'h1f == rd ? _next_reg_T_392 : _GEN_4421; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:{46,46}]
  wire [63:0] _GEN_4462 = _T_783 ? _GEN_4423 : _GEN_4391; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4463 = _T_783 ? _GEN_4424 : _GEN_4392; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4464 = _T_783 ? _GEN_4425 : _GEN_4393; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4465 = _T_783 ? _GEN_4426 : _GEN_4394; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4466 = _T_783 ? _GEN_4427 : _GEN_4395; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4467 = _T_783 ? _GEN_4428 : _GEN_4396; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4468 = _T_783 ? _GEN_4429 : _GEN_4397; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4469 = _T_783 ? _GEN_4430 : _GEN_4398; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4470 = _T_783 ? _GEN_4431 : _GEN_4399; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4471 = _T_783 ? _GEN_4432 : _GEN_4400; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4472 = _T_783 ? _GEN_4433 : _GEN_4401; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4473 = _T_783 ? _GEN_4434 : _GEN_4402; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4474 = _T_783 ? _GEN_4435 : _GEN_4403; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4475 = _T_783 ? _GEN_4436 : _GEN_4404; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4476 = _T_783 ? _GEN_4437 : _GEN_4405; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4477 = _T_783 ? _GEN_4438 : _GEN_4406; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4478 = _T_783 ? _GEN_4439 : _GEN_4407; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4479 = _T_783 ? _GEN_4440 : _GEN_4408; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4480 = _T_783 ? _GEN_4441 : _GEN_4409; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4481 = _T_783 ? _GEN_4442 : _GEN_4410; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4482 = _T_783 ? _GEN_4443 : _GEN_4411; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4483 = _T_783 ? _GEN_4444 : _GEN_4412; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4484 = _T_783 ? _GEN_4445 : _GEN_4413; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4485 = _T_783 ? _GEN_4446 : _GEN_4414; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4486 = _T_783 ? _GEN_4447 : _GEN_4415; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4487 = _T_783 ? _GEN_4448 : _GEN_4416; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4488 = _T_783 ? _GEN_4449 : _GEN_4417; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4489 = _T_783 ? _GEN_4450 : _GEN_4418; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4490 = _T_783 ? _GEN_4451 : _GEN_4419; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4491 = _T_783 ? _GEN_4452 : _GEN_4420; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [63:0] _GEN_4492 = _T_783 ? _GEN_4453 : _GEN_4421; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 398:22]
  wire [62:0] _GEN_5 = {{31'd0}, _GEN_101[31:0]}; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:78]
  wire [62:0] _next_reg_T_395 = _GEN_5 << _GEN_910[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:78]
  wire  next_reg_signBit_8 = _next_reg_T_395[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_398 = next_reg_signBit_8 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_399 = {_next_reg_T_398,_next_reg_T_395[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_4494 = 5'h1 == rd ? _next_reg_T_399 : _GEN_4462; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4495 = 5'h2 == rd ? _next_reg_T_399 : _GEN_4463; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4496 = 5'h3 == rd ? _next_reg_T_399 : _GEN_4464; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4497 = 5'h4 == rd ? _next_reg_T_399 : _GEN_4465; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4498 = 5'h5 == rd ? _next_reg_T_399 : _GEN_4466; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4499 = 5'h6 == rd ? _next_reg_T_399 : _GEN_4467; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4500 = 5'h7 == rd ? _next_reg_T_399 : _GEN_4468; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4501 = 5'h8 == rd ? _next_reg_T_399 : _GEN_4469; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4502 = 5'h9 == rd ? _next_reg_T_399 : _GEN_4470; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4503 = 5'ha == rd ? _next_reg_T_399 : _GEN_4471; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4504 = 5'hb == rd ? _next_reg_T_399 : _GEN_4472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4505 = 5'hc == rd ? _next_reg_T_399 : _GEN_4473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4506 = 5'hd == rd ? _next_reg_T_399 : _GEN_4474; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4507 = 5'he == rd ? _next_reg_T_399 : _GEN_4475; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4508 = 5'hf == rd ? _next_reg_T_399 : _GEN_4476; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4509 = 5'h10 == rd ? _next_reg_T_399 : _GEN_4477; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4510 = 5'h11 == rd ? _next_reg_T_399 : _GEN_4478; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4511 = 5'h12 == rd ? _next_reg_T_399 : _GEN_4479; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4512 = 5'h13 == rd ? _next_reg_T_399 : _GEN_4480; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4513 = 5'h14 == rd ? _next_reg_T_399 : _GEN_4481; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4514 = 5'h15 == rd ? _next_reg_T_399 : _GEN_4482; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4515 = 5'h16 == rd ? _next_reg_T_399 : _GEN_4483; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4516 = 5'h17 == rd ? _next_reg_T_399 : _GEN_4484; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4517 = 5'h18 == rd ? _next_reg_T_399 : _GEN_4485; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4518 = 5'h19 == rd ? _next_reg_T_399 : _GEN_4486; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4519 = 5'h1a == rd ? _next_reg_T_399 : _GEN_4487; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4520 = 5'h1b == rd ? _next_reg_T_399 : _GEN_4488; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4521 = 5'h1c == rd ? _next_reg_T_399 : _GEN_4489; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4522 = 5'h1d == rd ? _next_reg_T_399 : _GEN_4490; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4523 = 5'h1e == rd ? _next_reg_T_399 : _GEN_4491; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4524 = 5'h1f == rd ? _next_reg_T_399 : _GEN_4492; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:{46,46}]
  wire [63:0] _GEN_4533 = _T_790 ? _GEN_4494 : _GEN_4462; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4534 = _T_790 ? _GEN_4495 : _GEN_4463; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4535 = _T_790 ? _GEN_4496 : _GEN_4464; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4536 = _T_790 ? _GEN_4497 : _GEN_4465; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4537 = _T_790 ? _GEN_4498 : _GEN_4466; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4538 = _T_790 ? _GEN_4499 : _GEN_4467; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4539 = _T_790 ? _GEN_4500 : _GEN_4468; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4540 = _T_790 ? _GEN_4501 : _GEN_4469; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4541 = _T_790 ? _GEN_4502 : _GEN_4470; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4542 = _T_790 ? _GEN_4503 : _GEN_4471; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4543 = _T_790 ? _GEN_4504 : _GEN_4472; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4544 = _T_790 ? _GEN_4505 : _GEN_4473; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4545 = _T_790 ? _GEN_4506 : _GEN_4474; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4546 = _T_790 ? _GEN_4507 : _GEN_4475; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4547 = _T_790 ? _GEN_4508 : _GEN_4476; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4548 = _T_790 ? _GEN_4509 : _GEN_4477; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4549 = _T_790 ? _GEN_4510 : _GEN_4478; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4550 = _T_790 ? _GEN_4511 : _GEN_4479; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4551 = _T_790 ? _GEN_4512 : _GEN_4480; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4552 = _T_790 ? _GEN_4513 : _GEN_4481; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4553 = _T_790 ? _GEN_4514 : _GEN_4482; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4554 = _T_790 ? _GEN_4515 : _GEN_4483; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4555 = _T_790 ? _GEN_4516 : _GEN_4484; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4556 = _T_790 ? _GEN_4517 : _GEN_4485; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4557 = _T_790 ? _GEN_4518 : _GEN_4486; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4558 = _T_790 ? _GEN_4519 : _GEN_4487; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4559 = _T_790 ? _GEN_4520 : _GEN_4488; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4560 = _T_790 ? _GEN_4521 : _GEN_4489; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4561 = _T_790 ? _GEN_4522 : _GEN_4490; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4562 = _T_790 ? _GEN_4523 : _GEN_4491; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [63:0] _GEN_4563 = _T_790 ? _GEN_4524 : _GEN_4492; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 400:22]
  wire [31:0] _next_reg_T_402 = _GEN_101[31:0] >> _GEN_910[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:78]
  wire  next_reg_signBit_9 = _next_reg_T_402[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_405 = next_reg_signBit_9 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_406 = {_next_reg_T_405,_next_reg_T_402}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_4565 = 5'h1 == rd ? _next_reg_T_406 : _GEN_4533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4566 = 5'h2 == rd ? _next_reg_T_406 : _GEN_4534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4567 = 5'h3 == rd ? _next_reg_T_406 : _GEN_4535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4568 = 5'h4 == rd ? _next_reg_T_406 : _GEN_4536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4569 = 5'h5 == rd ? _next_reg_T_406 : _GEN_4537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4570 = 5'h6 == rd ? _next_reg_T_406 : _GEN_4538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4571 = 5'h7 == rd ? _next_reg_T_406 : _GEN_4539; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4572 = 5'h8 == rd ? _next_reg_T_406 : _GEN_4540; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4573 = 5'h9 == rd ? _next_reg_T_406 : _GEN_4541; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4574 = 5'ha == rd ? _next_reg_T_406 : _GEN_4542; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4575 = 5'hb == rd ? _next_reg_T_406 : _GEN_4543; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4576 = 5'hc == rd ? _next_reg_T_406 : _GEN_4544; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4577 = 5'hd == rd ? _next_reg_T_406 : _GEN_4545; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4578 = 5'he == rd ? _next_reg_T_406 : _GEN_4546; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4579 = 5'hf == rd ? _next_reg_T_406 : _GEN_4547; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4580 = 5'h10 == rd ? _next_reg_T_406 : _GEN_4548; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4581 = 5'h11 == rd ? _next_reg_T_406 : _GEN_4549; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4582 = 5'h12 == rd ? _next_reg_T_406 : _GEN_4550; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4583 = 5'h13 == rd ? _next_reg_T_406 : _GEN_4551; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4584 = 5'h14 == rd ? _next_reg_T_406 : _GEN_4552; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4585 = 5'h15 == rd ? _next_reg_T_406 : _GEN_4553; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4586 = 5'h16 == rd ? _next_reg_T_406 : _GEN_4554; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4587 = 5'h17 == rd ? _next_reg_T_406 : _GEN_4555; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4588 = 5'h18 == rd ? _next_reg_T_406 : _GEN_4556; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4589 = 5'h19 == rd ? _next_reg_T_406 : _GEN_4557; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4590 = 5'h1a == rd ? _next_reg_T_406 : _GEN_4558; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4591 = 5'h1b == rd ? _next_reg_T_406 : _GEN_4559; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4592 = 5'h1c == rd ? _next_reg_T_406 : _GEN_4560; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4593 = 5'h1d == rd ? _next_reg_T_406 : _GEN_4561; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4594 = 5'h1e == rd ? _next_reg_T_406 : _GEN_4562; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4595 = 5'h1f == rd ? _next_reg_T_406 : _GEN_4563; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:{46,46}]
  wire [63:0] _GEN_4604 = _T_797 ? _GEN_4565 : _GEN_4533; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4605 = _T_797 ? _GEN_4566 : _GEN_4534; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4606 = _T_797 ? _GEN_4567 : _GEN_4535; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4607 = _T_797 ? _GEN_4568 : _GEN_4536; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4608 = _T_797 ? _GEN_4569 : _GEN_4537; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4609 = _T_797 ? _GEN_4570 : _GEN_4538; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4610 = _T_797 ? _GEN_4571 : _GEN_4539; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4611 = _T_797 ? _GEN_4572 : _GEN_4540; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4612 = _T_797 ? _GEN_4573 : _GEN_4541; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4613 = _T_797 ? _GEN_4574 : _GEN_4542; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4614 = _T_797 ? _GEN_4575 : _GEN_4543; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4615 = _T_797 ? _GEN_4576 : _GEN_4544; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4616 = _T_797 ? _GEN_4577 : _GEN_4545; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4617 = _T_797 ? _GEN_4578 : _GEN_4546; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4618 = _T_797 ? _GEN_4579 : _GEN_4547; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4619 = _T_797 ? _GEN_4580 : _GEN_4548; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4620 = _T_797 ? _GEN_4581 : _GEN_4549; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4621 = _T_797 ? _GEN_4582 : _GEN_4550; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4622 = _T_797 ? _GEN_4583 : _GEN_4551; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4623 = _T_797 ? _GEN_4584 : _GEN_4552; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4624 = _T_797 ? _GEN_4585 : _GEN_4553; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4625 = _T_797 ? _GEN_4586 : _GEN_4554; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4626 = _T_797 ? _GEN_4587 : _GEN_4555; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4627 = _T_797 ? _GEN_4588 : _GEN_4556; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4628 = _T_797 ? _GEN_4589 : _GEN_4557; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4629 = _T_797 ? _GEN_4590 : _GEN_4558; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4630 = _T_797 ? _GEN_4591 : _GEN_4559; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4631 = _T_797 ? _GEN_4592 : _GEN_4560; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4632 = _T_797 ? _GEN_4593 : _GEN_4561; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4633 = _T_797 ? _GEN_4594 : _GEN_4562; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [63:0] _GEN_4634 = _T_797 ? _GEN_4595 : _GEN_4563; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 401:22]
  wire [31:0] _next_reg_T_410 = _GEN_101[31:0] - _GEN_910[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:78]
  wire  next_reg_signBit_10 = _next_reg_T_410[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_413 = next_reg_signBit_10 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_414 = {_next_reg_T_413,_next_reg_T_410}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_4636 = 5'h1 == rd ? _next_reg_T_414 : _GEN_4604; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4637 = 5'h2 == rd ? _next_reg_T_414 : _GEN_4605; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4638 = 5'h3 == rd ? _next_reg_T_414 : _GEN_4606; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4639 = 5'h4 == rd ? _next_reg_T_414 : _GEN_4607; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4640 = 5'h5 == rd ? _next_reg_T_414 : _GEN_4608; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4641 = 5'h6 == rd ? _next_reg_T_414 : _GEN_4609; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4642 = 5'h7 == rd ? _next_reg_T_414 : _GEN_4610; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4643 = 5'h8 == rd ? _next_reg_T_414 : _GEN_4611; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4644 = 5'h9 == rd ? _next_reg_T_414 : _GEN_4612; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4645 = 5'ha == rd ? _next_reg_T_414 : _GEN_4613; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4646 = 5'hb == rd ? _next_reg_T_414 : _GEN_4614; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4647 = 5'hc == rd ? _next_reg_T_414 : _GEN_4615; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4648 = 5'hd == rd ? _next_reg_T_414 : _GEN_4616; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4649 = 5'he == rd ? _next_reg_T_414 : _GEN_4617; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4650 = 5'hf == rd ? _next_reg_T_414 : _GEN_4618; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4651 = 5'h10 == rd ? _next_reg_T_414 : _GEN_4619; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4652 = 5'h11 == rd ? _next_reg_T_414 : _GEN_4620; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4653 = 5'h12 == rd ? _next_reg_T_414 : _GEN_4621; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4654 = 5'h13 == rd ? _next_reg_T_414 : _GEN_4622; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4655 = 5'h14 == rd ? _next_reg_T_414 : _GEN_4623; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4656 = 5'h15 == rd ? _next_reg_T_414 : _GEN_4624; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4657 = 5'h16 == rd ? _next_reg_T_414 : _GEN_4625; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4658 = 5'h17 == rd ? _next_reg_T_414 : _GEN_4626; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4659 = 5'h18 == rd ? _next_reg_T_414 : _GEN_4627; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4660 = 5'h19 == rd ? _next_reg_T_414 : _GEN_4628; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4661 = 5'h1a == rd ? _next_reg_T_414 : _GEN_4629; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4662 = 5'h1b == rd ? _next_reg_T_414 : _GEN_4630; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4663 = 5'h1c == rd ? _next_reg_T_414 : _GEN_4631; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4664 = 5'h1d == rd ? _next_reg_T_414 : _GEN_4632; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4665 = 5'h1e == rd ? _next_reg_T_414 : _GEN_4633; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4666 = 5'h1f == rd ? _next_reg_T_414 : _GEN_4634; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:{46,46}]
  wire [63:0] _GEN_4675 = _T_804 ? _GEN_4636 : _GEN_4604; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4676 = _T_804 ? _GEN_4637 : _GEN_4605; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4677 = _T_804 ? _GEN_4638 : _GEN_4606; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4678 = _T_804 ? _GEN_4639 : _GEN_4607; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4679 = _T_804 ? _GEN_4640 : _GEN_4608; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4680 = _T_804 ? _GEN_4641 : _GEN_4609; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4681 = _T_804 ? _GEN_4642 : _GEN_4610; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4682 = _T_804 ? _GEN_4643 : _GEN_4611; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4683 = _T_804 ? _GEN_4644 : _GEN_4612; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4684 = _T_804 ? _GEN_4645 : _GEN_4613; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4685 = _T_804 ? _GEN_4646 : _GEN_4614; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4686 = _T_804 ? _GEN_4647 : _GEN_4615; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4687 = _T_804 ? _GEN_4648 : _GEN_4616; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4688 = _T_804 ? _GEN_4649 : _GEN_4617; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4689 = _T_804 ? _GEN_4650 : _GEN_4618; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4690 = _T_804 ? _GEN_4651 : _GEN_4619; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4691 = _T_804 ? _GEN_4652 : _GEN_4620; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4692 = _T_804 ? _GEN_4653 : _GEN_4621; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4693 = _T_804 ? _GEN_4654 : _GEN_4622; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4694 = _T_804 ? _GEN_4655 : _GEN_4623; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4695 = _T_804 ? _GEN_4656 : _GEN_4624; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4696 = _T_804 ? _GEN_4657 : _GEN_4625; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4697 = _T_804 ? _GEN_4658 : _GEN_4626; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4698 = _T_804 ? _GEN_4659 : _GEN_4627; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4699 = _T_804 ? _GEN_4660 : _GEN_4628; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4700 = _T_804 ? _GEN_4661 : _GEN_4629; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4701 = _T_804 ? _GEN_4662 : _GEN_4630; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4702 = _T_804 ? _GEN_4663 : _GEN_4631; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4703 = _T_804 ? _GEN_4664 : _GEN_4632; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4704 = _T_804 ? _GEN_4665 : _GEN_4633; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [63:0] _GEN_4705 = _T_804 ? _GEN_4666 : _GEN_4634; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 403:22]
  wire [31:0] _next_reg_T_419 = $signed(_next_reg_T_370) >>> _GEN_910[4:0]; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:108]
  wire  next_reg_signBit_11 = _next_reg_T_419[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_421 = next_reg_signBit_11 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_422 = {_next_reg_T_421,_next_reg_T_419}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_4707 = 5'h1 == rd ? _next_reg_T_422 : _GEN_4675; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4708 = 5'h2 == rd ? _next_reg_T_422 : _GEN_4676; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4709 = 5'h3 == rd ? _next_reg_T_422 : _GEN_4677; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4710 = 5'h4 == rd ? _next_reg_T_422 : _GEN_4678; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4711 = 5'h5 == rd ? _next_reg_T_422 : _GEN_4679; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4712 = 5'h6 == rd ? _next_reg_T_422 : _GEN_4680; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4713 = 5'h7 == rd ? _next_reg_T_422 : _GEN_4681; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4714 = 5'h8 == rd ? _next_reg_T_422 : _GEN_4682; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4715 = 5'h9 == rd ? _next_reg_T_422 : _GEN_4683; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4716 = 5'ha == rd ? _next_reg_T_422 : _GEN_4684; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4717 = 5'hb == rd ? _next_reg_T_422 : _GEN_4685; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4718 = 5'hc == rd ? _next_reg_T_422 : _GEN_4686; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4719 = 5'hd == rd ? _next_reg_T_422 : _GEN_4687; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4720 = 5'he == rd ? _next_reg_T_422 : _GEN_4688; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4721 = 5'hf == rd ? _next_reg_T_422 : _GEN_4689; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4722 = 5'h10 == rd ? _next_reg_T_422 : _GEN_4690; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4723 = 5'h11 == rd ? _next_reg_T_422 : _GEN_4691; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4724 = 5'h12 == rd ? _next_reg_T_422 : _GEN_4692; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4725 = 5'h13 == rd ? _next_reg_T_422 : _GEN_4693; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4726 = 5'h14 == rd ? _next_reg_T_422 : _GEN_4694; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4727 = 5'h15 == rd ? _next_reg_T_422 : _GEN_4695; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4728 = 5'h16 == rd ? _next_reg_T_422 : _GEN_4696; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4729 = 5'h17 == rd ? _next_reg_T_422 : _GEN_4697; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4730 = 5'h18 == rd ? _next_reg_T_422 : _GEN_4698; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4731 = 5'h19 == rd ? _next_reg_T_422 : _GEN_4699; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4732 = 5'h1a == rd ? _next_reg_T_422 : _GEN_4700; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4733 = 5'h1b == rd ? _next_reg_T_422 : _GEN_4701; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4734 = 5'h1c == rd ? _next_reg_T_422 : _GEN_4702; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4735 = 5'h1d == rd ? _next_reg_T_422 : _GEN_4703; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4736 = 5'h1e == rd ? _next_reg_T_422 : _GEN_4704; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4737 = 5'h1f == rd ? _next_reg_T_422 : _GEN_4705; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:{46,46}]
  wire [63:0] _GEN_4746 = _T_811 ? _GEN_4707 : _GEN_4675; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4747 = _T_811 ? _GEN_4708 : _GEN_4676; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4748 = _T_811 ? _GEN_4709 : _GEN_4677; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4749 = _T_811 ? _GEN_4710 : _GEN_4678; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4750 = _T_811 ? _GEN_4711 : _GEN_4679; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4751 = _T_811 ? _GEN_4712 : _GEN_4680; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4752 = _T_811 ? _GEN_4713 : _GEN_4681; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4753 = _T_811 ? _GEN_4714 : _GEN_4682; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4754 = _T_811 ? _GEN_4715 : _GEN_4683; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4755 = _T_811 ? _GEN_4716 : _GEN_4684; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4756 = _T_811 ? _GEN_4717 : _GEN_4685; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4757 = _T_811 ? _GEN_4718 : _GEN_4686; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4758 = _T_811 ? _GEN_4719 : _GEN_4687; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4759 = _T_811 ? _GEN_4720 : _GEN_4688; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4760 = _T_811 ? _GEN_4721 : _GEN_4689; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4761 = _T_811 ? _GEN_4722 : _GEN_4690; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4762 = _T_811 ? _GEN_4723 : _GEN_4691; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4763 = _T_811 ? _GEN_4724 : _GEN_4692; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4764 = _T_811 ? _GEN_4725 : _GEN_4693; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4765 = _T_811 ? _GEN_4726 : _GEN_4694; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4766 = _T_811 ? _GEN_4727 : _GEN_4695; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4767 = _T_811 ? _GEN_4728 : _GEN_4696; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4768 = _T_811 ? _GEN_4729 : _GEN_4697; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4769 = _T_811 ? _GEN_4730 : _GEN_4698; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4770 = _T_811 ? _GEN_4731 : _GEN_4699; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4771 = _T_811 ? _GEN_4732 : _GEN_4700; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4772 = _T_811 ? _GEN_4733 : _GEN_4701; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4773 = _T_811 ? _GEN_4734 : _GEN_4702; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4774 = _T_811 ? _GEN_4735 : _GEN_4703; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4775 = _T_811 ? _GEN_4736 : _GEN_4704; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire [63:0] _GEN_4776 = _T_811 ? _GEN_4737 : _GEN_4705; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 404:22]
  wire  _GEN_4800 = next_reg_LevelVec_10_1_valid | _GEN_3660; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_4801 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec__1_addr : _GEN_3661; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire  _GEN_4811 = next_reg_LevelVec_10_0_valid | _GEN_3663; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_4812 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec__0_addr : _GEN_3664; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] _GEN_4870 = next_reg_success_10 ? next_reg_finaladdr : _GEN_3177; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 69:25]
  wire  _GEN_4872 = next_reg_success_10 ? _GEN_3702 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_4873 = next_reg_vmEnable_10 | _GEN_3657; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_4874 = next_reg_vmEnable_10 ? next_reg_LevelVec__2_addr : _GEN_3658; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_4876 = next_reg_vmEnable_10 ? _GEN_4800 : _GEN_3660; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_4877 = next_reg_vmEnable_10 ? _GEN_4801 : _GEN_3661; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_4879 = next_reg_vmEnable_10 ? _GEN_4811 : _GEN_3663; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_4880 = next_reg_vmEnable_10 ? _GEN_4812 : _GEN_3664; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_4886 = next_reg_vmEnable_10 ? _GEN_4870 : _T_844; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22 74:23]
  wire  _GEN_4888 = next_reg_vmEnable_10 ? _GEN_4872 : _GEN_3702; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _next_reg_T_480 = {32'h0,_next_reg_T_221[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [63:0] _GEN_4890 = 5'h1 == rd ? _next_reg_T_480 : _GEN_4746; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4891 = 5'h2 == rd ? _next_reg_T_480 : _GEN_4747; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4892 = 5'h3 == rd ? _next_reg_T_480 : _GEN_4748; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4893 = 5'h4 == rd ? _next_reg_T_480 : _GEN_4749; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4894 = 5'h5 == rd ? _next_reg_T_480 : _GEN_4750; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4895 = 5'h6 == rd ? _next_reg_T_480 : _GEN_4751; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4896 = 5'h7 == rd ? _next_reg_T_480 : _GEN_4752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4897 = 5'h8 == rd ? _next_reg_T_480 : _GEN_4753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4898 = 5'h9 == rd ? _next_reg_T_480 : _GEN_4754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4899 = 5'ha == rd ? _next_reg_T_480 : _GEN_4755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4900 = 5'hb == rd ? _next_reg_T_480 : _GEN_4756; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4901 = 5'hc == rd ? _next_reg_T_480 : _GEN_4757; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4902 = 5'hd == rd ? _next_reg_T_480 : _GEN_4758; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4903 = 5'he == rd ? _next_reg_T_480 : _GEN_4759; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4904 = 5'hf == rd ? _next_reg_T_480 : _GEN_4760; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4905 = 5'h10 == rd ? _next_reg_T_480 : _GEN_4761; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4906 = 5'h11 == rd ? _next_reg_T_480 : _GEN_4762; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4907 = 5'h12 == rd ? _next_reg_T_480 : _GEN_4763; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4908 = 5'h13 == rd ? _next_reg_T_480 : _GEN_4764; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4909 = 5'h14 == rd ? _next_reg_T_480 : _GEN_4765; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4910 = 5'h15 == rd ? _next_reg_T_480 : _GEN_4766; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4911 = 5'h16 == rd ? _next_reg_T_480 : _GEN_4767; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4912 = 5'h17 == rd ? _next_reg_T_480 : _GEN_4768; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4913 = 5'h18 == rd ? _next_reg_T_480 : _GEN_4769; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4914 = 5'h19 == rd ? _next_reg_T_480 : _GEN_4770; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4915 = 5'h1a == rd ? _next_reg_T_480 : _GEN_4771; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4916 = 5'h1b == rd ? _next_reg_T_480 : _GEN_4772; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4917 = 5'h1c == rd ? _next_reg_T_480 : _GEN_4773; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4918 = 5'h1d == rd ? _next_reg_T_480 : _GEN_4774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4919 = 5'h1e == rd ? _next_reg_T_480 : _GEN_4775; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire [63:0] _GEN_4920 = 5'h1f == rd ? _next_reg_T_480 : _GEN_4776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 412:{22,22}]
  wire  _GEN_4921 = _T_848 | _GEN_3163; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 63:22]
  wire  _GEN_4922 = _T_848 ? _GEN_4873 : _GEN_3657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4923 = _T_848 ? _GEN_4874 : _GEN_3658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire  _GEN_4925 = _T_848 ? _GEN_4876 : _GEN_3660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4926 = _T_848 ? _GEN_4877 : _GEN_3661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire  _GEN_4928 = _T_848 ? _GEN_4879 : _GEN_3663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4929 = _T_848 ? _GEN_4880 : _GEN_3664; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4935 = _T_848 ? _GEN_4886 : _T_844; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55 414:23]
  wire  _GEN_4937 = _T_848 ? _GEN_4888 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [6:0] _GEN_4938 = _T_848 ? 7'h20 : _GEN_3180; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 76:25]
  wire [63:0] _GEN_4940 = _T_848 ? _GEN_4890 : _GEN_4746; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4941 = _T_848 ? _GEN_4891 : _GEN_4747; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4942 = _T_848 ? _GEN_4892 : _GEN_4748; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4943 = _T_848 ? _GEN_4893 : _GEN_4749; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4944 = _T_848 ? _GEN_4894 : _GEN_4750; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4945 = _T_848 ? _GEN_4895 : _GEN_4751; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4946 = _T_848 ? _GEN_4896 : _GEN_4752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4947 = _T_848 ? _GEN_4897 : _GEN_4753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4948 = _T_848 ? _GEN_4898 : _GEN_4754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4949 = _T_848 ? _GEN_4899 : _GEN_4755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4950 = _T_848 ? _GEN_4900 : _GEN_4756; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4951 = _T_848 ? _GEN_4901 : _GEN_4757; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4952 = _T_848 ? _GEN_4902 : _GEN_4758; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4953 = _T_848 ? _GEN_4903 : _GEN_4759; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4954 = _T_848 ? _GEN_4904 : _GEN_4760; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4955 = _T_848 ? _GEN_4905 : _GEN_4761; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4956 = _T_848 ? _GEN_4906 : _GEN_4762; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4957 = _T_848 ? _GEN_4907 : _GEN_4763; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4958 = _T_848 ? _GEN_4908 : _GEN_4764; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4959 = _T_848 ? _GEN_4909 : _GEN_4765; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4960 = _T_848 ? _GEN_4910 : _GEN_4766; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4961 = _T_848 ? _GEN_4911 : _GEN_4767; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4962 = _T_848 ? _GEN_4912 : _GEN_4768; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4963 = _T_848 ? _GEN_4913 : _GEN_4769; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4964 = _T_848 ? _GEN_4914 : _GEN_4770; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4965 = _T_848 ? _GEN_4915 : _GEN_4771; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4966 = _T_848 ? _GEN_4916 : _GEN_4772; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4967 = _T_848 ? _GEN_4917 : _GEN_4773; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4968 = _T_848 ? _GEN_4918 : _GEN_4774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4969 = _T_848 ? _GEN_4919 : _GEN_4775; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire [63:0] _GEN_4970 = _T_848 ? _GEN_4920 : _GEN_4776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 411:55]
  wire  _GEN_4979 = _T_818 ? _GEN_4921 : _GEN_3163; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire  _GEN_4980 = _T_818 ? _GEN_4922 : _GEN_3657; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_4981 = _T_818 ? _GEN_4923 : _GEN_3658; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire  _GEN_4983 = _T_818 ? _GEN_4925 : _GEN_3660; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_4984 = _T_818 ? _GEN_4926 : _GEN_3661; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire  _GEN_4986 = _T_818 ? _GEN_4928 : _GEN_3663; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_4987 = _T_818 ? _GEN_4929 : _GEN_3664; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_4993 = _T_818 ? _GEN_4935 : _GEN_3177; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire  _GEN_4995 = _T_818 ? _GEN_4937 : _GEN_3702; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [6:0] _GEN_4996 = _T_818 ? _GEN_4938 : _GEN_3180; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_4998 = _T_818 ? _GEN_4940 : _GEN_4746; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_4999 = _T_818 ? _GEN_4941 : _GEN_4747; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5000 = _T_818 ? _GEN_4942 : _GEN_4748; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5001 = _T_818 ? _GEN_4943 : _GEN_4749; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5002 = _T_818 ? _GEN_4944 : _GEN_4750; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5003 = _T_818 ? _GEN_4945 : _GEN_4751; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5004 = _T_818 ? _GEN_4946 : _GEN_4752; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5005 = _T_818 ? _GEN_4947 : _GEN_4753; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5006 = _T_818 ? _GEN_4948 : _GEN_4754; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5007 = _T_818 ? _GEN_4949 : _GEN_4755; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5008 = _T_818 ? _GEN_4950 : _GEN_4756; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5009 = _T_818 ? _GEN_4951 : _GEN_4757; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5010 = _T_818 ? _GEN_4952 : _GEN_4758; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5011 = _T_818 ? _GEN_4953 : _GEN_4759; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5012 = _T_818 ? _GEN_4954 : _GEN_4760; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5013 = _T_818 ? _GEN_4955 : _GEN_4761; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5014 = _T_818 ? _GEN_4956 : _GEN_4762; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5015 = _T_818 ? _GEN_4957 : _GEN_4763; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5016 = _T_818 ? _GEN_4958 : _GEN_4764; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5017 = _T_818 ? _GEN_4959 : _GEN_4765; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5018 = _T_818 ? _GEN_4960 : _GEN_4766; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5019 = _T_818 ? _GEN_4961 : _GEN_4767; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5020 = _T_818 ? _GEN_4962 : _GEN_4768; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5021 = _T_818 ? _GEN_4963 : _GEN_4769; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5022 = _T_818 ? _GEN_4964 : _GEN_4770; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5023 = _T_818 ? _GEN_4965 : _GEN_4771; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5024 = _T_818 ? _GEN_4966 : _GEN_4772; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5025 = _T_818 ? _GEN_4967 : _GEN_4773; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5026 = _T_818 ? _GEN_4968 : _GEN_4774; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5027 = _T_818 ? _GEN_4969 : _GEN_4775; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire [63:0] _GEN_5028 = _T_818 ? _GEN_4970 : _GEN_4776; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 409:21]
  wire  _GEN_5053 = next_reg_LevelVec_10_1_valid | _GEN_4983; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_5054 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec__1_addr : _GEN_4984; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire  _GEN_5064 = next_reg_LevelVec_10_0_valid | _GEN_4986; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_5065 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec__0_addr : _GEN_4987; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] _GEN_5123 = next_reg_success_10 ? next_reg_finaladdr : _GEN_4993; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 69:25]
  wire  _GEN_5125 = next_reg_success_10 ? _GEN_4995 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5126 = next_reg_vmEnable_10 | _GEN_4980; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_5127 = next_reg_vmEnable_10 ? next_reg_LevelVec__2_addr : _GEN_4981; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_5129 = next_reg_vmEnable_10 ? _GEN_5053 : _GEN_4983; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_5130 = next_reg_vmEnable_10 ? _GEN_5054 : _GEN_4984; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_5132 = next_reg_vmEnable_10 ? _GEN_5064 : _GEN_4986; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_5133 = next_reg_vmEnable_10 ? _GEN_5065 : _GEN_4987; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_5139 = next_reg_vmEnable_10 ? _GEN_5123 : _T_844; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22 74:23]
  wire  _GEN_5141 = next_reg_vmEnable_10 ? _GEN_5125 : _GEN_4995; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_5143 = 5'h1 == rd ? _next_reg_T_100 : _GEN_4998; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5144 = 5'h2 == rd ? _next_reg_T_100 : _GEN_4999; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5145 = 5'h3 == rd ? _next_reg_T_100 : _GEN_5000; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5146 = 5'h4 == rd ? _next_reg_T_100 : _GEN_5001; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5147 = 5'h5 == rd ? _next_reg_T_100 : _GEN_5002; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5148 = 5'h6 == rd ? _next_reg_T_100 : _GEN_5003; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5149 = 5'h7 == rd ? _next_reg_T_100 : _GEN_5004; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5150 = 5'h8 == rd ? _next_reg_T_100 : _GEN_5005; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5151 = 5'h9 == rd ? _next_reg_T_100 : _GEN_5006; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5152 = 5'ha == rd ? _next_reg_T_100 : _GEN_5007; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5153 = 5'hb == rd ? _next_reg_T_100 : _GEN_5008; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5154 = 5'hc == rd ? _next_reg_T_100 : _GEN_5009; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5155 = 5'hd == rd ? _next_reg_T_100 : _GEN_5010; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5156 = 5'he == rd ? _next_reg_T_100 : _GEN_5011; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5157 = 5'hf == rd ? _next_reg_T_100 : _GEN_5012; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5158 = 5'h10 == rd ? _next_reg_T_100 : _GEN_5013; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5159 = 5'h11 == rd ? _next_reg_T_100 : _GEN_5014; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5160 = 5'h12 == rd ? _next_reg_T_100 : _GEN_5015; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5161 = 5'h13 == rd ? _next_reg_T_100 : _GEN_5016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5162 = 5'h14 == rd ? _next_reg_T_100 : _GEN_5017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5163 = 5'h15 == rd ? _next_reg_T_100 : _GEN_5018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5164 = 5'h16 == rd ? _next_reg_T_100 : _GEN_5019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5165 = 5'h17 == rd ? _next_reg_T_100 : _GEN_5020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5166 = 5'h18 == rd ? _next_reg_T_100 : _GEN_5021; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5167 = 5'h19 == rd ? _next_reg_T_100 : _GEN_5022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5168 = 5'h1a == rd ? _next_reg_T_100 : _GEN_5023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5169 = 5'h1b == rd ? _next_reg_T_100 : _GEN_5024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5170 = 5'h1c == rd ? _next_reg_T_100 : _GEN_5025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5171 = 5'h1d == rd ? _next_reg_T_100 : _GEN_5026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5172 = 5'h1e == rd ? _next_reg_T_100 : _GEN_5027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire [63:0] _GEN_5173 = 5'h1f == rd ? _next_reg_T_100 : _GEN_5028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 421:{22,22}]
  wire  _GEN_5174 = _T_850 | _GEN_4979; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 63:22]
  wire  _GEN_5175 = _T_850 ? _GEN_5126 : _GEN_4980; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5176 = _T_850 ? _GEN_5127 : _GEN_4981; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire  _GEN_5178 = _T_850 ? _GEN_5129 : _GEN_4983; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5179 = _T_850 ? _GEN_5130 : _GEN_4984; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire  _GEN_5181 = _T_850 ? _GEN_5132 : _GEN_4986; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5182 = _T_850 ? _GEN_5133 : _GEN_4987; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5188 = _T_850 ? _GEN_5139 : _T_844; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55 423:23]
  wire  _GEN_5190 = _T_850 ? _GEN_5141 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [6:0] _GEN_5191 = _T_850 ? 7'h40 : _GEN_4996; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 76:25]
  wire [63:0] _GEN_5193 = _T_850 ? _GEN_5143 : _GEN_4998; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5194 = _T_850 ? _GEN_5144 : _GEN_4999; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5195 = _T_850 ? _GEN_5145 : _GEN_5000; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5196 = _T_850 ? _GEN_5146 : _GEN_5001; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5197 = _T_850 ? _GEN_5147 : _GEN_5002; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5198 = _T_850 ? _GEN_5148 : _GEN_5003; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5199 = _T_850 ? _GEN_5149 : _GEN_5004; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5200 = _T_850 ? _GEN_5150 : _GEN_5005; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5201 = _T_850 ? _GEN_5151 : _GEN_5006; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5202 = _T_850 ? _GEN_5152 : _GEN_5007; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5203 = _T_850 ? _GEN_5153 : _GEN_5008; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5204 = _T_850 ? _GEN_5154 : _GEN_5009; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5205 = _T_850 ? _GEN_5155 : _GEN_5010; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5206 = _T_850 ? _GEN_5156 : _GEN_5011; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5207 = _T_850 ? _GEN_5157 : _GEN_5012; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5208 = _T_850 ? _GEN_5158 : _GEN_5013; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5209 = _T_850 ? _GEN_5159 : _GEN_5014; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5210 = _T_850 ? _GEN_5160 : _GEN_5015; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5211 = _T_850 ? _GEN_5161 : _GEN_5016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5212 = _T_850 ? _GEN_5162 : _GEN_5017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5213 = _T_850 ? _GEN_5163 : _GEN_5018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5214 = _T_850 ? _GEN_5164 : _GEN_5019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5215 = _T_850 ? _GEN_5165 : _GEN_5020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5216 = _T_850 ? _GEN_5166 : _GEN_5021; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5217 = _T_850 ? _GEN_5167 : _GEN_5022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5218 = _T_850 ? _GEN_5168 : _GEN_5023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5219 = _T_850 ? _GEN_5169 : _GEN_5024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5220 = _T_850 ? _GEN_5170 : _GEN_5025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5221 = _T_850 ? _GEN_5171 : _GEN_5026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5222 = _T_850 ? _GEN_5172 : _GEN_5027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire [63:0] _GEN_5223 = _T_850 ? _GEN_5173 : _GEN_5028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 420:55]
  wire  _GEN_5232 = _T_838 ? _GEN_5174 : _GEN_4979; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire  _GEN_5233 = _T_838 ? _GEN_5175 : _GEN_4980; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5234 = _T_838 ? _GEN_5176 : _GEN_4981; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire  _GEN_5236 = _T_838 ? _GEN_5178 : _GEN_4983; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5237 = _T_838 ? _GEN_5179 : _GEN_4984; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire  _GEN_5239 = _T_838 ? _GEN_5181 : _GEN_4986; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5240 = _T_838 ? _GEN_5182 : _GEN_4987; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5246 = _T_838 ? _GEN_5188 : _GEN_4993; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire  _GEN_5248 = _T_838 ? _GEN_5190 : _GEN_4995; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [6:0] _GEN_5249 = _T_838 ? _GEN_5191 : _GEN_4996; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5251 = _T_838 ? _GEN_5193 : _GEN_4998; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5252 = _T_838 ? _GEN_5194 : _GEN_4999; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5253 = _T_838 ? _GEN_5195 : _GEN_5000; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5254 = _T_838 ? _GEN_5196 : _GEN_5001; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5255 = _T_838 ? _GEN_5197 : _GEN_5002; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5256 = _T_838 ? _GEN_5198 : _GEN_5003; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5257 = _T_838 ? _GEN_5199 : _GEN_5004; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5258 = _T_838 ? _GEN_5200 : _GEN_5005; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5259 = _T_838 ? _GEN_5201 : _GEN_5006; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5260 = _T_838 ? _GEN_5202 : _GEN_5007; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5261 = _T_838 ? _GEN_5203 : _GEN_5008; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5262 = _T_838 ? _GEN_5204 : _GEN_5009; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5263 = _T_838 ? _GEN_5205 : _GEN_5010; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5264 = _T_838 ? _GEN_5206 : _GEN_5011; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5265 = _T_838 ? _GEN_5207 : _GEN_5012; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5266 = _T_838 ? _GEN_5208 : _GEN_5013; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5267 = _T_838 ? _GEN_5209 : _GEN_5014; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5268 = _T_838 ? _GEN_5210 : _GEN_5015; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5269 = _T_838 ? _GEN_5211 : _GEN_5016; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5270 = _T_838 ? _GEN_5212 : _GEN_5017; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5271 = _T_838 ? _GEN_5213 : _GEN_5018; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5272 = _T_838 ? _GEN_5214 : _GEN_5019; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5273 = _T_838 ? _GEN_5215 : _GEN_5020; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5274 = _T_838 ? _GEN_5216 : _GEN_5021; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5275 = _T_838 ? _GEN_5217 : _GEN_5022; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5276 = _T_838 ? _GEN_5218 : _GEN_5023; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5277 = _T_838 ? _GEN_5219 : _GEN_5024; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5278 = _T_838 ? _GEN_5220 : _GEN_5025; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5279 = _T_838 ? _GEN_5221 : _GEN_5026; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5280 = _T_838 ? _GEN_5222 : _GEN_5027; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire [63:0] _GEN_5281 = _T_838 ? _GEN_5223 : _GEN_5028; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 418:20]
  wire  _GEN_5306 = next_reg_LevelVec_10_1_valid | _GEN_5236; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_5307 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec__1_addr : _GEN_5237; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire  _GEN_5317 = next_reg_LevelVec_10_0_valid | _GEN_5239; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_5318 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec__0_addr : _GEN_5240; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] _GEN_5376 = success_8 ? finaladdr_1 : _GEN_3670; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 97:26]
  wire  _GEN_5378 = success_8 ? _GEN_5248 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5379 = next_reg_vmEnable_10 | _GEN_5233; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_5380 = next_reg_vmEnable_10 ? next_reg_LevelVec__2_addr : _GEN_5234; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_5382 = next_reg_vmEnable_10 ? _GEN_5306 : _GEN_5236; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_5383 = next_reg_vmEnable_10 ? _GEN_5307 : _GEN_5237; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_5385 = next_reg_vmEnable_10 ? _GEN_5317 : _GEN_5239; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_5386 = next_reg_vmEnable_10 ? _GEN_5318 : _GEN_5240; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_5392 = next_reg_vmEnable_10 ? _GEN_5376 : _T_844; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22 102:24]
  wire  _GEN_5394 = next_reg_vmEnable_10 ? _GEN_5378 : _GEN_5248; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_5395 = _T_850 | _GEN_3656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 92:23]
  wire  _GEN_5396 = _T_850 ? _GEN_5379 : _GEN_5233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55]
  wire [63:0] _GEN_5397 = _T_850 ? _GEN_5380 : _GEN_5234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55]
  wire  _GEN_5399 = _T_850 ? _GEN_5382 : _GEN_5236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55]
  wire [63:0] _GEN_5400 = _T_850 ? _GEN_5383 : _GEN_5237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55]
  wire  _GEN_5402 = _T_850 ? _GEN_5385 : _GEN_5239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55]
  wire [63:0] _GEN_5403 = _T_850 ? _GEN_5386 : _GEN_5240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55]
  wire [63:0] _GEN_5409 = _T_850 ? _GEN_5392 : _T_844; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55 433:24]
  wire  _GEN_5411 = _T_850 ? _GEN_5394 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire [6:0] _GEN_5412 = _T_850 ? 7'h40 : _GEN_3673; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 104:26]
  wire [63:0] _GEN_5413 = _T_850 ? _GEN_910 : _GEN_3674; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 430:55 src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:26]
  wire  _GEN_5423 = _T_858 ? _GEN_5395 : _GEN_3656; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire  _GEN_5424 = _T_858 ? _GEN_5396 : _GEN_5233; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire [63:0] _GEN_5425 = _T_858 ? _GEN_5397 : _GEN_5234; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire  _GEN_5427 = _T_858 ? _GEN_5399 : _GEN_5236; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire [63:0] _GEN_5428 = _T_858 ? _GEN_5400 : _GEN_5237; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire  _GEN_5430 = _T_858 ? _GEN_5402 : _GEN_5239; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire [63:0] _GEN_5431 = _T_858 ? _GEN_5403 : _GEN_5240; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire [63:0] _GEN_5437 = _T_858 ? _GEN_5409 : _GEN_3670; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire  _GEN_5439 = _T_858 ? _GEN_5411 : _GEN_5248; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire [6:0] _GEN_5440 = _T_858 ? _GEN_5412 : _GEN_3673; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire [63:0] _GEN_5441 = _T_858 ? _GEN_5413 : _GEN_3674; // @[src/main/scala/rvspeccore/core/spec/instset/IBase.scala 428:20]
  wire [63:0] _next_reg_T_540 = io_now_reg_2 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:52]
  wire [5:0] next_reg_rOff_7 = {_next_reg_T_540[2:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 58:51]
  wire [63:0] next_reg_LevelVec_7_2_addr = {8'h0,io_now_csr_satp[43:0],_next_reg_T_540[38:30],3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 268:31]
  wire [63:0] _next_reg_LevelVec_1_addr_T_31 = {8'h0,next_reg_PTE_30_ppn,_next_reg_T_540[29:21],3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 302:54]
  wire [63:0] _GEN_5444 = next_reg_PTEFlag_30_r | next_reg_PTEFlag_30_x ? 64'h0 : _next_reg_LevelVec_1_addr_T_31; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 287:42 292:47 302:48]
  wire [63:0] next_reg_LevelVec_7_1_addr = ~next_reg_PTEFlag_30_v | ~next_reg_PTEFlag_30_r & next_reg_PTEFlag_30_w ? 64'h0
     : _GEN_5444; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 277:57 282:45]
  wire [63:0] _next_reg_LevelVec_0_addr_T_31 = {8'h0,next_reg_PTE_31_ppn,_next_reg_T_540[20:12],3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 305:54]
  wire [63:0] _GEN_5459 = next_reg_PTEFlag_31_r | next_reg_PTEFlag_31_x ? 64'h0 : _next_reg_LevelVec_0_addr_T_31; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 287:42 292:47 305:48]
  wire [63:0] _GEN_5463 = ~next_reg_PTEFlag_31_v | ~next_reg_PTEFlag_31_r & next_reg_PTEFlag_31_w ? 64'h0 : _GEN_5459; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 277:57 282:45]
  wire  _GEN_5466 = next_reg_LevelVec_10_1_valid | _GEN_5427; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_5467 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec_7_1_addr : _GEN_5428; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] next_reg_LevelVec_7_0_addr = next_reg_LevelVec_10_1_valid ? _GEN_5463 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 271:41 317:43]
  wire  _GEN_5477 = next_reg_LevelVec_10_0_valid | _GEN_5430; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_5478 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec_7_0_addr : _GEN_5431; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [55:0] _next_reg_finaladdr_T_75 = {_GEN_8145[53:10],_next_reg_T_540[11:0]}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 364:31]
  wire [55:0] _next_reg_finaladdr_T_77 = _next_reg_finaladdr_T_75 & _GEN_11189; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 364:103]
  wire [63:0] _next_reg_finaladdr_T_78 = _next_reg_T_540 & _GEN_11190; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 366:26]
  wire [63:0] _GEN_11224 = {{8'd0}, _next_reg_finaladdr_T_77}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 366:18]
  wire [63:0] _next_reg_finaladdr_T_79 = _GEN_11224 | _next_reg_finaladdr_T_78; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 366:18]
  wire [63:0] _GEN_5504 = _next_reg_T_797 ? 64'h0 : _next_reg_finaladdr_T_79; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 349:99 352:26 364:23]
  wire [63:0] _GEN_5510 = next_reg_permLoad_10 ? _GEN_5504 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 346:11 372:24]
  wire [63:0] next_reg_finaladdr_7 = ~(next_reg_successLevel_10 == 2'h3) ? _GEN_5510 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 335:37 377:22]
  wire [63:0] _GEN_5536 = next_reg_success_10 ? next_reg_finaladdr_7 : _GEN_5246; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 69:25]
  wire  _GEN_5538 = next_reg_success_10 ? _GEN_5439 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5539 = next_reg_vmEnable_10 | _GEN_5424; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_5540 = next_reg_vmEnable_10 ? next_reg_LevelVec_7_2_addr : _GEN_5425; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_5542 = next_reg_vmEnable_10 ? _GEN_5466 : _GEN_5427; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_5543 = next_reg_vmEnable_10 ? _GEN_5467 : _GEN_5428; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_5545 = next_reg_vmEnable_10 ? _GEN_5477 : _GEN_5430; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_5546 = next_reg_vmEnable_10 ? _GEN_5478 : _GEN_5431; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_5552 = next_reg_vmEnable_10 ? _GEN_5536 : _next_reg_T_540; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22 74:23]
  wire  _GEN_5554 = next_reg_vmEnable_10 ? _GEN_5538 : _GEN_5439; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _next_reg_T_593 = io_mem_read_data >> next_reg_rOff_7; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 77:22]
  wire [63:0] _next_reg_T_594 = _next_reg_T_593 & 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 77:31]
  wire  next_reg_signBit_13 = _next_reg_T_594[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_597 = next_reg_signBit_13 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_598 = {_next_reg_T_597,_next_reg_T_594[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_5556 = 5'h1 == rd ? _next_reg_T_598 : _GEN_5251; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5557 = 5'h2 == rd ? _next_reg_T_598 : _GEN_5252; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5558 = 5'h3 == rd ? _next_reg_T_598 : _GEN_5253; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5559 = 5'h4 == rd ? _next_reg_T_598 : _GEN_5254; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5560 = 5'h5 == rd ? _next_reg_T_598 : _GEN_5255; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5561 = 5'h6 == rd ? _next_reg_T_598 : _GEN_5256; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5562 = 5'h7 == rd ? _next_reg_T_598 : _GEN_5257; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5563 = 5'h8 == rd ? _next_reg_T_598 : _GEN_5258; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5564 = 5'h9 == rd ? _next_reg_T_598 : _GEN_5259; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5565 = 5'ha == rd ? _next_reg_T_598 : _GEN_5260; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5566 = 5'hb == rd ? _next_reg_T_598 : _GEN_5261; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5567 = 5'hc == rd ? _next_reg_T_598 : _GEN_5262; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5568 = 5'hd == rd ? _next_reg_T_598 : _GEN_5263; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5569 = 5'he == rd ? _next_reg_T_598 : _GEN_5264; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5570 = 5'hf == rd ? _next_reg_T_598 : _GEN_5265; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5571 = 5'h10 == rd ? _next_reg_T_598 : _GEN_5266; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5572 = 5'h11 == rd ? _next_reg_T_598 : _GEN_5267; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5573 = 5'h12 == rd ? _next_reg_T_598 : _GEN_5268; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5574 = 5'h13 == rd ? _next_reg_T_598 : _GEN_5269; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5575 = 5'h14 == rd ? _next_reg_T_598 : _GEN_5270; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5576 = 5'h15 == rd ? _next_reg_T_598 : _GEN_5271; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5577 = 5'h16 == rd ? _next_reg_T_598 : _GEN_5272; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5578 = 5'h17 == rd ? _next_reg_T_598 : _GEN_5273; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5579 = 5'h18 == rd ? _next_reg_T_598 : _GEN_5274; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5580 = 5'h19 == rd ? _next_reg_T_598 : _GEN_5275; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5581 = 5'h1a == rd ? _next_reg_T_598 : _GEN_5276; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5582 = 5'h1b == rd ? _next_reg_T_598 : _GEN_5277; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5583 = 5'h1c == rd ? _next_reg_T_598 : _GEN_5278; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5584 = 5'h1d == rd ? _next_reg_T_598 : _GEN_5279; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5585 = 5'h1e == rd ? _next_reg_T_598 : _GEN_5280; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire [63:0] _GEN_5586 = 5'h1f == rd ? _next_reg_T_598 : _GEN_5281; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 141:{20,20}]
  wire  _GEN_5595 = _T_937 | _GEN_5232; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 63:22]
  wire  _GEN_5596 = _T_937 ? _GEN_5539 : _GEN_5424; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5597 = _T_937 ? _GEN_5540 : _GEN_5425; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire  _GEN_5599 = _T_937 ? _GEN_5542 : _GEN_5427; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5600 = _T_937 ? _GEN_5543 : _GEN_5428; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire  _GEN_5602 = _T_937 ? _GEN_5545 : _GEN_5430; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5603 = _T_937 ? _GEN_5546 : _GEN_5431; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5609 = _T_937 ? _GEN_5552 : _GEN_5246; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire  _GEN_5611 = _T_937 ? _GEN_5554 : _GEN_5439; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [6:0] _GEN_5612 = _T_937 ? 7'h20 : _GEN_5249; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 76:25]
  wire [63:0] _GEN_5614 = _T_937 ? _GEN_5556 : _GEN_5251; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5615 = _T_937 ? _GEN_5557 : _GEN_5252; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5616 = _T_937 ? _GEN_5558 : _GEN_5253; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5617 = _T_937 ? _GEN_5559 : _GEN_5254; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5618 = _T_937 ? _GEN_5560 : _GEN_5255; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5619 = _T_937 ? _GEN_5561 : _GEN_5256; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5620 = _T_937 ? _GEN_5562 : _GEN_5257; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5621 = _T_937 ? _GEN_5563 : _GEN_5258; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5622 = _T_937 ? _GEN_5564 : _GEN_5259; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5623 = _T_937 ? _GEN_5565 : _GEN_5260; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5624 = _T_937 ? _GEN_5566 : _GEN_5261; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5625 = _T_937 ? _GEN_5567 : _GEN_5262; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5626 = _T_937 ? _GEN_5568 : _GEN_5263; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5627 = _T_937 ? _GEN_5569 : _GEN_5264; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5628 = _T_937 ? _GEN_5570 : _GEN_5265; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5629 = _T_937 ? _GEN_5571 : _GEN_5266; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5630 = _T_937 ? _GEN_5572 : _GEN_5267; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5631 = _T_937 ? _GEN_5573 : _GEN_5268; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5632 = _T_937 ? _GEN_5574 : _GEN_5269; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5633 = _T_937 ? _GEN_5575 : _GEN_5270; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5634 = _T_937 ? _GEN_5576 : _GEN_5271; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5635 = _T_937 ? _GEN_5577 : _GEN_5272; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5636 = _T_937 ? _GEN_5578 : _GEN_5273; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5637 = _T_937 ? _GEN_5579 : _GEN_5274; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5638 = _T_937 ? _GEN_5580 : _GEN_5275; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5639 = _T_937 ? _GEN_5581 : _GEN_5276; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5640 = _T_937 ? _GEN_5582 : _GEN_5277; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5641 = _T_937 ? _GEN_5583 : _GEN_5278; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5642 = _T_937 ? _GEN_5584 : _GEN_5279; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5643 = _T_937 ? _GEN_5585 : _GEN_5280; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire [63:0] _GEN_5644 = _T_937 ? _GEN_5586 : _GEN_5281; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 138:24]
  wire  _GEN_5668 = next_reg_LevelVec_10_1_valid | _GEN_5599; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_5669 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec_7_1_addr : _GEN_5600; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire  _GEN_5679 = next_reg_LevelVec_10_0_valid | _GEN_5602; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_5680 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec_7_0_addr : _GEN_5603; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] _GEN_5712 = next_reg_permStore_10 ? _GEN_5504 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 346:11 372:24]
  wire [63:0] finaladdr_5 = ~(next_reg_successLevel_10 == 2'h3) ? _GEN_5712 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 335:37 377:22]
  wire [63:0] _GEN_5738 = success_8 ? finaladdr_5 : _GEN_5437; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 97:26]
  wire  _GEN_5740 = success_8 ? _GEN_5611 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5741 = next_reg_vmEnable_10 | _GEN_5596; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_5742 = next_reg_vmEnable_10 ? next_reg_LevelVec_7_2_addr : _GEN_5597; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_5744 = next_reg_vmEnable_10 ? _GEN_5668 : _GEN_5599; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_5745 = next_reg_vmEnable_10 ? _GEN_5669 : _GEN_5600; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_5747 = next_reg_vmEnable_10 ? _GEN_5679 : _GEN_5602; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_5748 = next_reg_vmEnable_10 ? _GEN_5680 : _GEN_5603; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_5754 = next_reg_vmEnable_10 ? _GEN_5738 : _next_reg_T_540; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22 102:24]
  wire  _GEN_5756 = next_reg_vmEnable_10 ? _GEN_5740 : _GEN_5611; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_5763 = _T_944 | _GEN_5423; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 92:23]
  wire  _GEN_5764 = _T_944 ? _GEN_5741 : _GEN_5596; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24]
  wire [63:0] _GEN_5765 = _T_944 ? _GEN_5742 : _GEN_5597; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24]
  wire  _GEN_5767 = _T_944 ? _GEN_5744 : _GEN_5599; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24]
  wire [63:0] _GEN_5768 = _T_944 ? _GEN_5745 : _GEN_5600; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24]
  wire  _GEN_5770 = _T_944 ? _GEN_5747 : _GEN_5602; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24]
  wire [63:0] _GEN_5771 = _T_944 ? _GEN_5748 : _GEN_5603; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24]
  wire [63:0] _GEN_5777 = _T_944 ? _GEN_5754 : _GEN_5437; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24]
  wire  _GEN_5779 = _T_944 ? _GEN_5756 : _GEN_5611; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24]
  wire [6:0] _GEN_5780 = _T_944 ? 7'h20 : _GEN_5440; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 104:26]
  wire [63:0] _GEN_5781 = _T_944 ? {{32'd0}, _GEN_910[31:0]} : _GEN_5441; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 143:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:26]
  wire [2:0] _GEN_5961 = _T_1005 ? inst[9:7] : 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 99:24]
  wire [2:0] _GEN_6195 = _T_1014 ? inst[9:7] : _GEN_5961; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_6288 = _T_1107 ? inst[9:7] : _GEN_6195; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_6332 = _T_1116 ? inst[9:7] : _GEN_6288; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_6801 = _T_1212 ? inst[9:7] : _GEN_6332; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_6905 = _T_1226 ? inst[9:7] : _GEN_6801; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_7009 = _T_1234 ? inst[9:7] : _GEN_6905; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_7284 = _T_1266 ? inst[9:7] : _GEN_7009; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_7419 = _T_1274 ? inst[9:7] : _GEN_7284; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_7554 = _T_1282 ? inst[9:7] : _GEN_7419; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_7689 = _T_1290 ? inst[9:7] : _GEN_7554; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_8251 = _T_1376 ? inst[9:7] : _GEN_7689; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_8485 = _T_1385 ? inst[9:7] : _GEN_8251; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_8679 = _T_1459 ? inst[9:7] : _GEN_8485; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_8814 = _T_1467 ? inst[9:7] : _GEN_8679; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] rs1P = io_valid ? _GEN_8814 : 3'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 99:24]
  wire [2:0] _GEN_5963 = _T_1005 ? inst[4:2] : 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 98:24]
  wire [2:0] _GEN_6291 = _T_1107 ? rs1P : _GEN_5963; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:111 186:24]
  wire [2:0] _GEN_6335 = _T_1116 ? rs1P : _GEN_6291; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:111 194:24]
  wire [2:0] _GEN_6628 = _T_1183 ? inst[4:2] : _GEN_6335; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_6804 = _T_1212 ? rs1P : _GEN_6628; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:111 235:24]
  wire [2:0] _GEN_6908 = _T_1226 ? rs1P : _GEN_6804; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:111 240:24]
  wire [2:0] _GEN_7012 = _T_1234 ? rs1P : _GEN_6908; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 119:111 245:24]
  wire [2:0] _GEN_7288 = _T_1266 ? rs1P : _GEN_7012; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:111 253:23]
  wire [2:0] _GEN_7423 = _T_1274 ? rs1P : _GEN_7288; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:111 254:23]
  wire [2:0] _GEN_7558 = _T_1282 ? rs1P : _GEN_7423; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:111 255:23]
  wire [2:0] _GEN_7693 = _T_1290 ? rs1P : _GEN_7558; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:111 256:23]
  wire [2:0] _GEN_8253 = _T_1376 ? inst[4:2] : _GEN_7693; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_8683 = _T_1459 ? rs1P : _GEN_8253; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:111 297:24]
  wire [2:0] _GEN_8818 = _T_1467 ? rs1P : _GEN_8683; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 118:111 301:24]
  wire [2:0] rdP = io_valid ? _GEN_8818 : 3'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 98:24]
  wire [4:0] _T_1012 = {2'h1,rdP}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [4:0] _next_reg_T_599 = {2'h1,rs1P}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire [63:0] _GEN_5783 = 5'h1 == _next_reg_T_599 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5784 = 5'h2 == _next_reg_T_599 ? io_now_reg_2 : _GEN_5783; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5785 = 5'h3 == _next_reg_T_599 ? io_now_reg_3 : _GEN_5784; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5786 = 5'h4 == _next_reg_T_599 ? io_now_reg_4 : _GEN_5785; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5787 = 5'h5 == _next_reg_T_599 ? io_now_reg_5 : _GEN_5786; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5788 = 5'h6 == _next_reg_T_599 ? io_now_reg_6 : _GEN_5787; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5789 = 5'h7 == _next_reg_T_599 ? io_now_reg_7 : _GEN_5788; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5790 = 5'h8 == _next_reg_T_599 ? io_now_reg_8 : _GEN_5789; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5791 = 5'h9 == _next_reg_T_599 ? io_now_reg_9 : _GEN_5790; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5792 = 5'ha == _next_reg_T_599 ? io_now_reg_10 : _GEN_5791; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5793 = 5'hb == _next_reg_T_599 ? io_now_reg_11 : _GEN_5792; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5794 = 5'hc == _next_reg_T_599 ? io_now_reg_12 : _GEN_5793; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5795 = 5'hd == _next_reg_T_599 ? io_now_reg_13 : _GEN_5794; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5796 = 5'he == _next_reg_T_599 ? io_now_reg_14 : _GEN_5795; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5797 = 5'hf == _next_reg_T_599 ? io_now_reg_15 : _GEN_5796; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5798 = 5'h10 == _next_reg_T_599 ? io_now_reg_16 : _GEN_5797; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5799 = 5'h11 == _next_reg_T_599 ? io_now_reg_17 : _GEN_5798; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5800 = 5'h12 == _next_reg_T_599 ? io_now_reg_18 : _GEN_5799; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5801 = 5'h13 == _next_reg_T_599 ? io_now_reg_19 : _GEN_5800; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5802 = 5'h14 == _next_reg_T_599 ? io_now_reg_20 : _GEN_5801; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5803 = 5'h15 == _next_reg_T_599 ? io_now_reg_21 : _GEN_5802; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5804 = 5'h16 == _next_reg_T_599 ? io_now_reg_22 : _GEN_5803; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5805 = 5'h17 == _next_reg_T_599 ? io_now_reg_23 : _GEN_5804; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5806 = 5'h18 == _next_reg_T_599 ? io_now_reg_24 : _GEN_5805; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5807 = 5'h19 == _next_reg_T_599 ? io_now_reg_25 : _GEN_5806; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5808 = 5'h1a == _next_reg_T_599 ? io_now_reg_26 : _GEN_5807; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5809 = 5'h1b == _next_reg_T_599 ? io_now_reg_27 : _GEN_5808; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5810 = 5'h1c == _next_reg_T_599 ? io_now_reg_28 : _GEN_5809; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5811 = 5'h1d == _next_reg_T_599 ? io_now_reg_29 : _GEN_5810; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5812 = 5'h1e == _next_reg_T_599 ? io_now_reg_30 : _GEN_5811; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _GEN_5813 = 5'h1f == _next_reg_T_599 ? io_now_reg_31 : _GEN_5812; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{68,68}]
  wire [63:0] _next_reg_T_601 = _GEN_5813 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:68]
  wire [5:0] next_reg_rOff_8 = {_next_reg_T_601[2:0], 3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 58:51]
  wire [63:0] next_reg_LevelVec_8_2_addr = {8'h0,io_now_csr_satp[43:0],_next_reg_T_601[38:30],3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 268:31]
  wire [63:0] _next_reg_LevelVec_1_addr_T_35 = {8'h0,next_reg_PTE_30_ppn,_next_reg_T_601[29:21],3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 302:54]
  wire [63:0] _GEN_5815 = next_reg_PTEFlag_30_r | next_reg_PTEFlag_30_x ? 64'h0 : _next_reg_LevelVec_1_addr_T_35; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 287:42 292:47 302:48]
  wire [63:0] next_reg_LevelVec_8_1_addr = ~next_reg_PTEFlag_30_v | ~next_reg_PTEFlag_30_r & next_reg_PTEFlag_30_w ? 64'h0
     : _GEN_5815; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 277:57 282:45]
  wire [63:0] _next_reg_LevelVec_0_addr_T_35 = {8'h0,next_reg_PTE_31_ppn,_next_reg_T_601[20:12],3'h0}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 305:54]
  wire [63:0] _GEN_5830 = next_reg_PTEFlag_31_r | next_reg_PTEFlag_31_x ? 64'h0 : _next_reg_LevelVec_0_addr_T_35; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 287:42 292:47 305:48]
  wire [63:0] _GEN_5834 = ~next_reg_PTEFlag_31_v | ~next_reg_PTEFlag_31_r & next_reg_PTEFlag_31_w ? 64'h0 : _GEN_5830; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 277:57 282:45]
  wire  _GEN_5837 = next_reg_LevelVec_10_1_valid | _GEN_5767; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_5838 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec_8_1_addr : _GEN_5768; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] next_reg_LevelVec_8_0_addr = next_reg_LevelVec_10_1_valid ? _GEN_5834 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 271:41 317:43]
  wire  _GEN_5848 = next_reg_LevelVec_10_0_valid | _GEN_5770; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_5849 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec_8_0_addr : _GEN_5771; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [55:0] _next_reg_finaladdr_T_85 = {_GEN_8145[53:10],_next_reg_T_601[11:0]}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 364:31]
  wire [55:0] _next_reg_finaladdr_T_87 = _next_reg_finaladdr_T_85 & _GEN_11189; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 364:103]
  wire [63:0] _next_reg_finaladdr_T_88 = _next_reg_T_601 & _GEN_11190; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 366:26]
  wire [63:0] _GEN_11230 = {{8'd0}, _next_reg_finaladdr_T_87}; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 366:18]
  wire [63:0] _next_reg_finaladdr_T_89 = _GEN_11230 | _next_reg_finaladdr_T_88; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 366:18]
  wire [63:0] _GEN_5875 = _next_reg_T_797 ? 64'h0 : _next_reg_finaladdr_T_89; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 349:99 352:26 364:23]
  wire [63:0] _GEN_5881 = next_reg_permLoad_10 ? _GEN_5875 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 346:11 372:24]
  wire [63:0] next_reg_finaladdr_8 = ~(next_reg_successLevel_10 == 2'h3) ? _GEN_5881 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 335:37 377:22]
  wire [63:0] _GEN_5907 = next_reg_success_10 ? next_reg_finaladdr_8 : _GEN_5609; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 69:25]
  wire  _GEN_5909 = next_reg_success_10 ? _GEN_5779 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_5910 = next_reg_vmEnable_10 | _GEN_5764; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_5911 = next_reg_vmEnable_10 ? next_reg_LevelVec_8_2_addr : _GEN_5765; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_5913 = next_reg_vmEnable_10 ? _GEN_5837 : _GEN_5767; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_5914 = next_reg_vmEnable_10 ? _GEN_5838 : _GEN_5768; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_5916 = next_reg_vmEnable_10 ? _GEN_5848 : _GEN_5770; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_5917 = next_reg_vmEnable_10 ? _GEN_5849 : _GEN_5771; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_5923 = next_reg_vmEnable_10 ? _GEN_5907 : _next_reg_T_601; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22 74:23]
  wire  _GEN_5925 = next_reg_vmEnable_10 ? _GEN_5909 : _GEN_5779; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _next_reg_T_654 = io_mem_read_data >> next_reg_rOff_8; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 77:22]
  wire [63:0] _next_reg_T_655 = _next_reg_T_654 & 64'hffffffff; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 77:31]
  wire  next_reg_signBit_14 = _next_reg_T_655[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_658 = next_reg_signBit_14 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_659 = {_next_reg_T_658,_next_reg_T_655[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_5927 = 5'h1 == _T_1012 ? _next_reg_T_659 : _GEN_5614; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5928 = 5'h2 == _T_1012 ? _next_reg_T_659 : _GEN_5615; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5929 = 5'h3 == _T_1012 ? _next_reg_T_659 : _GEN_5616; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5930 = 5'h4 == _T_1012 ? _next_reg_T_659 : _GEN_5617; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5931 = 5'h5 == _T_1012 ? _next_reg_T_659 : _GEN_5618; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5932 = 5'h6 == _T_1012 ? _next_reg_T_659 : _GEN_5619; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5933 = 5'h7 == _T_1012 ? _next_reg_T_659 : _GEN_5620; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5934 = 5'h8 == _T_1012 ? _next_reg_T_659 : _GEN_5621; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5935 = 5'h9 == _T_1012 ? _next_reg_T_659 : _GEN_5622; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5936 = 5'ha == _T_1012 ? _next_reg_T_659 : _GEN_5623; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5937 = 5'hb == _T_1012 ? _next_reg_T_659 : _GEN_5624; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5938 = 5'hc == _T_1012 ? _next_reg_T_659 : _GEN_5625; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5939 = 5'hd == _T_1012 ? _next_reg_T_659 : _GEN_5626; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5940 = 5'he == _T_1012 ? _next_reg_T_659 : _GEN_5627; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5941 = 5'hf == _T_1012 ? _next_reg_T_659 : _GEN_5628; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5942 = 5'h10 == _T_1012 ? _next_reg_T_659 : _GEN_5629; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5943 = 5'h11 == _T_1012 ? _next_reg_T_659 : _GEN_5630; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5944 = 5'h12 == _T_1012 ? _next_reg_T_659 : _GEN_5631; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5945 = 5'h13 == _T_1012 ? _next_reg_T_659 : _GEN_5632; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5946 = 5'h14 == _T_1012 ? _next_reg_T_659 : _GEN_5633; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5947 = 5'h15 == _T_1012 ? _next_reg_T_659 : _GEN_5634; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5948 = 5'h16 == _T_1012 ? _next_reg_T_659 : _GEN_5635; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5949 = 5'h17 == _T_1012 ? _next_reg_T_659 : _GEN_5636; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5950 = 5'h18 == _T_1012 ? _next_reg_T_659 : _GEN_5637; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5951 = 5'h19 == _T_1012 ? _next_reg_T_659 : _GEN_5638; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5952 = 5'h1a == _T_1012 ? _next_reg_T_659 : _GEN_5639; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5953 = 5'h1b == _T_1012 ? _next_reg_T_659 : _GEN_5640; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5954 = 5'h1c == _T_1012 ? _next_reg_T_659 : _GEN_5641; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5955 = 5'h1d == _T_1012 ? _next_reg_T_659 : _GEN_5642; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5956 = 5'h1e == _T_1012 ? _next_reg_T_659 : _GEN_5643; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire [63:0] _GEN_5957 = 5'h1f == _T_1012 ? _next_reg_T_659 : _GEN_5644; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 152:{28,28}]
  wire  _GEN_5966 = _T_1005 | _GEN_5595; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 63:22]
  wire  _GEN_5967 = _T_1005 ? _GEN_5910 : _GEN_5764; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5968 = _T_1005 ? _GEN_5911 : _GEN_5765; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire  _GEN_5970 = _T_1005 ? _GEN_5913 : _GEN_5767; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5971 = _T_1005 ? _GEN_5914 : _GEN_5768; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire  _GEN_5973 = _T_1005 ? _GEN_5916 : _GEN_5770; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5974 = _T_1005 ? _GEN_5917 : _GEN_5771; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5980 = _T_1005 ? _GEN_5923 : _GEN_5609; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire  _GEN_5982 = _T_1005 ? _GEN_5925 : _GEN_5779; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [6:0] _GEN_5983 = _T_1005 ? 7'h20 : _GEN_5612; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 76:25]
  wire [63:0] _GEN_5985 = _T_1005 ? _GEN_5927 : _GEN_5614; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5986 = _T_1005 ? _GEN_5928 : _GEN_5615; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5987 = _T_1005 ? _GEN_5929 : _GEN_5616; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5988 = _T_1005 ? _GEN_5930 : _GEN_5617; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5989 = _T_1005 ? _GEN_5931 : _GEN_5618; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5990 = _T_1005 ? _GEN_5932 : _GEN_5619; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5991 = _T_1005 ? _GEN_5933 : _GEN_5620; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5992 = _T_1005 ? _GEN_5934 : _GEN_5621; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5993 = _T_1005 ? _GEN_5935 : _GEN_5622; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5994 = _T_1005 ? _GEN_5936 : _GEN_5623; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5995 = _T_1005 ? _GEN_5937 : _GEN_5624; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5996 = _T_1005 ? _GEN_5938 : _GEN_5625; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5997 = _T_1005 ? _GEN_5939 : _GEN_5626; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5998 = _T_1005 ? _GEN_5940 : _GEN_5627; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_5999 = _T_1005 ? _GEN_5941 : _GEN_5628; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_6000 = _T_1005 ? _GEN_5942 : _GEN_5629; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_6001 = _T_1005 ? _GEN_5943 : _GEN_5630; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_6002 = _T_1005 ? _GEN_5944 : _GEN_5631; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_6003 = _T_1005 ? _GEN_5945 : _GEN_5632; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_6004 = _T_1005 ? _GEN_5946 : _GEN_5633; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_6005 = _T_1005 ? _GEN_5947 : _GEN_5634; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_6006 = _T_1005 ? _GEN_5948 : _GEN_5635; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_6007 = _T_1005 ? _GEN_5949 : _GEN_5636; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_6008 = _T_1005 ? _GEN_5950 : _GEN_5637; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_6009 = _T_1005 ? _GEN_5951 : _GEN_5638; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_6010 = _T_1005 ? _GEN_5952 : _GEN_5639; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_6011 = _T_1005 ? _GEN_5953 : _GEN_5640; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_6012 = _T_1005 ? _GEN_5954 : _GEN_5641; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_6013 = _T_1005 ? _GEN_5955 : _GEN_5642; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_6014 = _T_1005 ? _GEN_5956 : _GEN_5643; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [63:0] _GEN_6015 = _T_1005 ? _GEN_5957 : _GEN_5644; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 149:22]
  wire [2:0] _GEN_6197 = _T_1014 ? inst[4:2] : 3'h0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 100:24]
  wire [2:0] _GEN_7286 = _T_1266 ? inst[4:2] : _GEN_6197; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_7421 = _T_1274 ? inst[4:2] : _GEN_7286; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_7556 = _T_1282 ? inst[4:2] : _GEN_7421; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_7691 = _T_1290 ? inst[4:2] : _GEN_7556; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_8487 = _T_1385 ? inst[4:2] : _GEN_7691; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_8681 = _T_1459 ? inst[4:2] : _GEN_8487; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] _GEN_8816 = _T_1467 ? inst[4:2] : _GEN_8681; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24 src/main/scala/rvspeccore/core/tool/BitTool.scala 31:14]
  wire [2:0] rs2P = io_valid ? _GEN_8816 : 3'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 100:24]
  wire [4:0] _T_1024 = {2'h1,rs2P}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 133:33]
  wire  _GEN_6071 = next_reg_LevelVec_10_1_valid | _GEN_5970; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_6072 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec_8_1_addr : _GEN_5971; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire  _GEN_6082 = next_reg_LevelVec_10_0_valid | _GEN_5973; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_6083 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec_8_0_addr : _GEN_5974; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] _GEN_6115 = next_reg_permStore_10 ? _GEN_5875 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 346:11 372:24]
  wire [63:0] finaladdr_6 = ~(next_reg_successLevel_10 == 2'h3) ? _GEN_6115 : 64'h0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 335:37 377:22]
  wire [63:0] _GEN_6141 = success_8 ? finaladdr_6 : _GEN_5777; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 97:26]
  wire  _GEN_6143 = success_8 ? _GEN_5982 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_6144 = next_reg_vmEnable_10 | _GEN_5967; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_6145 = next_reg_vmEnable_10 ? next_reg_LevelVec_8_2_addr : _GEN_5968; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_6147 = next_reg_vmEnable_10 ? _GEN_6071 : _GEN_5970; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_6148 = next_reg_vmEnable_10 ? _GEN_6072 : _GEN_5971; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_6150 = next_reg_vmEnable_10 ? _GEN_6082 : _GEN_5973; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_6151 = next_reg_vmEnable_10 ? _GEN_6083 : _GEN_5974; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_6157 = next_reg_vmEnable_10 ? _GEN_6141 : _next_reg_T_601; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22 102:24]
  wire  _GEN_6159 = next_reg_vmEnable_10 ? _GEN_6143 : _GEN_5982; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_6161 = 5'h1 == _T_1024 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6162 = 5'h2 == _T_1024 ? io_now_reg_2 : _GEN_6161; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6163 = 5'h3 == _T_1024 ? io_now_reg_3 : _GEN_6162; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6164 = 5'h4 == _T_1024 ? io_now_reg_4 : _GEN_6163; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6165 = 5'h5 == _T_1024 ? io_now_reg_5 : _GEN_6164; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6166 = 5'h6 == _T_1024 ? io_now_reg_6 : _GEN_6165; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6167 = 5'h7 == _T_1024 ? io_now_reg_7 : _GEN_6166; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6168 = 5'h8 == _T_1024 ? io_now_reg_8 : _GEN_6167; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6169 = 5'h9 == _T_1024 ? io_now_reg_9 : _GEN_6168; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6170 = 5'ha == _T_1024 ? io_now_reg_10 : _GEN_6169; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6171 = 5'hb == _T_1024 ? io_now_reg_11 : _GEN_6170; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6172 = 5'hc == _T_1024 ? io_now_reg_12 : _GEN_6171; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6173 = 5'hd == _T_1024 ? io_now_reg_13 : _GEN_6172; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6174 = 5'he == _T_1024 ? io_now_reg_14 : _GEN_6173; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6175 = 5'hf == _T_1024 ? io_now_reg_15 : _GEN_6174; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6176 = 5'h10 == _T_1024 ? io_now_reg_16 : _GEN_6175; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6177 = 5'h11 == _T_1024 ? io_now_reg_17 : _GEN_6176; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6178 = 5'h12 == _T_1024 ? io_now_reg_18 : _GEN_6177; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6179 = 5'h13 == _T_1024 ? io_now_reg_19 : _GEN_6178; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6180 = 5'h14 == _T_1024 ? io_now_reg_20 : _GEN_6179; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6181 = 5'h15 == _T_1024 ? io_now_reg_21 : _GEN_6180; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6182 = 5'h16 == _T_1024 ? io_now_reg_22 : _GEN_6181; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6183 = 5'h17 == _T_1024 ? io_now_reg_23 : _GEN_6182; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6184 = 5'h18 == _T_1024 ? io_now_reg_24 : _GEN_6183; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6185 = 5'h19 == _T_1024 ? io_now_reg_25 : _GEN_6184; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6186 = 5'h1a == _T_1024 ? io_now_reg_26 : _GEN_6185; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6187 = 5'h1b == _T_1024 ? io_now_reg_27 : _GEN_6186; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6188 = 5'h1c == _T_1024 ? io_now_reg_28 : _GEN_6187; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6189 = 5'h1d == _T_1024 ? io_now_reg_29 : _GEN_6188; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6190 = 5'h1e == _T_1024 ? io_now_reg_30 : _GEN_6189; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire [63:0] _GEN_6191 = 5'h1f == _T_1024 ? io_now_reg_31 : _GEN_6190; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:{26,26}]
  wire  _GEN_6200 = _T_1014 | _GEN_5763; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 92:23]
  wire  _GEN_6201 = _T_1014 ? _GEN_6144 : _GEN_5967; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22]
  wire [63:0] _GEN_6202 = _T_1014 ? _GEN_6145 : _GEN_5968; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22]
  wire  _GEN_6204 = _T_1014 ? _GEN_6147 : _GEN_5970; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22]
  wire [63:0] _GEN_6205 = _T_1014 ? _GEN_6148 : _GEN_5971; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22]
  wire  _GEN_6207 = _T_1014 ? _GEN_6150 : _GEN_5973; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22]
  wire [63:0] _GEN_6208 = _T_1014 ? _GEN_6151 : _GEN_5974; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22]
  wire [63:0] _GEN_6214 = _T_1014 ? _GEN_6157 : _GEN_5777; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22]
  wire  _GEN_6216 = _T_1014 ? _GEN_6159 : _GEN_5982; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22]
  wire [6:0] _GEN_6217 = _T_1014 ? 7'h20 : _GEN_5780; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 104:26]
  wire [63:0] _GEN_6218 = _T_1014 ? _GEN_6191 : _GEN_5781; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 154:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:26]
  wire  _GEN_6224 = _T_1078 | _GEN_1993; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 160:21 163:25]
  wire [63:0] _GEN_6225 = _T_1078 ? _T_359 : _GEN_1994; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 160:21 164:25]
  wire [63:0] _next_reg_1_T_1 = io_now_pc + 64'h2; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 171:35]
  wire [63:0] _next_pc_T_23 = {_GEN_101[63:1],1'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 177:21]
  wire  _GEN_6240 = _T_1092 | _GEN_6224; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 175:25]
  wire [63:0] _GEN_6241 = _T_1092 ? _next_pc_T_23 : _GEN_6225; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 173:22 177:15]
  wire  _GEN_6248 = _T_1101 | _GEN_6240; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 181:25]
  wire [63:0] _GEN_6249 = _T_1101 ? _next_pc_T_23 : _GEN_6241; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 183:21]
  wire [63:0] _GEN_6250 = _T_1101 ? _next_reg_1_T_1 : _GEN_5985; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 179:24 184:21]
  wire  _GEN_6283 = _GEN_5813 == 64'h0 | _GEN_6248; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:42 190:27]
  wire [63:0] _GEN_6284 = _GEN_5813 == 64'h0 ? _T_359 : _GEN_6249; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 189:42 191:27]
  wire  _GEN_6293 = _T_1107 ? _GEN_6283 : _GEN_6248; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24]
  wire [63:0] _GEN_6294 = _T_1107 ? _GEN_6284 : _GEN_6249; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 186:24]
  wire  _GEN_6327 = _GEN_5813 != 64'h0 | _GEN_6293; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:42 198:27]
  wire [63:0] _GEN_6328 = _GEN_5813 != 64'h0 ? _T_359 : _GEN_6294; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 197:42 199:27]
  wire  _GEN_6337 = _T_1116 ? _GEN_6327 : _GEN_6293; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24]
  wire [63:0] _GEN_6338 = _T_1116 ? _GEN_6328 : _GEN_6294; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 194:24]
  wire [63:0] _GEN_6340 = 5'h1 == rd ? imm : _GEN_6250; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6341 = 5'h2 == rd ? imm : _GEN_5986; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6342 = 5'h3 == rd ? imm : _GEN_5987; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6343 = 5'h4 == rd ? imm : _GEN_5988; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6344 = 5'h5 == rd ? imm : _GEN_5989; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6345 = 5'h6 == rd ? imm : _GEN_5990; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6346 = 5'h7 == rd ? imm : _GEN_5991; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6347 = 5'h8 == rd ? imm : _GEN_5992; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6348 = 5'h9 == rd ? imm : _GEN_5993; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6349 = 5'ha == rd ? imm : _GEN_5994; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6350 = 5'hb == rd ? imm : _GEN_5995; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6351 = 5'hc == rd ? imm : _GEN_5996; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6352 = 5'hd == rd ? imm : _GEN_5997; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6353 = 5'he == rd ? imm : _GEN_5998; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6354 = 5'hf == rd ? imm : _GEN_5999; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6355 = 5'h10 == rd ? imm : _GEN_6000; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6356 = 5'h11 == rd ? imm : _GEN_6001; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6357 = 5'h12 == rd ? imm : _GEN_6002; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6358 = 5'h13 == rd ? imm : _GEN_6003; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6359 = 5'h14 == rd ? imm : _GEN_6004; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6360 = 5'h15 == rd ? imm : _GEN_6005; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6361 = 5'h16 == rd ? imm : _GEN_6006; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6362 = 5'h17 == rd ? imm : _GEN_6007; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6363 = 5'h18 == rd ? imm : _GEN_6008; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6364 = 5'h19 == rd ? imm : _GEN_6009; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6365 = 5'h1a == rd ? imm : _GEN_6010; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6366 = 5'h1b == rd ? imm : _GEN_6011; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6367 = 5'h1c == rd ? imm : _GEN_6012; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6368 = 5'h1d == rd ? imm : _GEN_6013; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6369 = 5'h1e == rd ? imm : _GEN_6014; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6370 = 5'h1f == rd ? imm : _GEN_6015; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 207:{20,20}]
  wire [63:0] _GEN_6380 = _T_1128 ? _GEN_6340 : _GEN_6250; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6381 = _T_1128 ? _GEN_6341 : _GEN_5986; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6382 = _T_1128 ? _GEN_6342 : _GEN_5987; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6383 = _T_1128 ? _GEN_6343 : _GEN_5988; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6384 = _T_1128 ? _GEN_6344 : _GEN_5989; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6385 = _T_1128 ? _GEN_6345 : _GEN_5990; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6386 = _T_1128 ? _GEN_6346 : _GEN_5991; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6387 = _T_1128 ? _GEN_6347 : _GEN_5992; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6388 = _T_1128 ? _GEN_6348 : _GEN_5993; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6389 = _T_1128 ? _GEN_6349 : _GEN_5994; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6390 = _T_1128 ? _GEN_6350 : _GEN_5995; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6391 = _T_1128 ? _GEN_6351 : _GEN_5996; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6392 = _T_1128 ? _GEN_6352 : _GEN_5997; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6393 = _T_1128 ? _GEN_6353 : _GEN_5998; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6394 = _T_1128 ? _GEN_6354 : _GEN_5999; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6395 = _T_1128 ? _GEN_6355 : _GEN_6000; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6396 = _T_1128 ? _GEN_6356 : _GEN_6001; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6397 = _T_1128 ? _GEN_6357 : _GEN_6002; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6398 = _T_1128 ? _GEN_6358 : _GEN_6003; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6399 = _T_1128 ? _GEN_6359 : _GEN_6004; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6400 = _T_1128 ? _GEN_6360 : _GEN_6005; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6401 = _T_1128 ? _GEN_6361 : _GEN_6006; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6402 = _T_1128 ? _GEN_6362 : _GEN_6007; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6403 = _T_1128 ? _GEN_6363 : _GEN_6008; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6404 = _T_1128 ? _GEN_6364 : _GEN_6009; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6405 = _T_1128 ? _GEN_6365 : _GEN_6010; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6406 = _T_1128 ? _GEN_6366 : _GEN_6011; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6407 = _T_1128 ? _GEN_6367 : _GEN_6012; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6408 = _T_1128 ? _GEN_6368 : _GEN_6013; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6409 = _T_1128 ? _GEN_6369 : _GEN_6014; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [63:0] _GEN_6410 = _T_1128 ? _GEN_6370 : _GEN_6015; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 204:22]
  wire [17:0] _nzimm_C_LUI_T_7 = {inst[12],inst[6],inst[5],inst[4],inst[3],inst[2],12'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire  nzimm_C_LUI_signBit = _nzimm_C_LUI_T_7[17]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [45:0] _nzimm_C_LUI_T_9 = nzimm_C_LUI_signBit ? 46'h3fffffffffff : 46'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] nzimm_C_LUI = {_nzimm_C_LUI_T_9,inst[12],inst[6],inst[5],inst[4],inst[3],inst[2],12'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_6412 = 5'h1 == rd ? nzimm_C_LUI : _GEN_6380; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6413 = 5'h2 == rd ? nzimm_C_LUI : _GEN_6381; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6414 = 5'h3 == rd ? nzimm_C_LUI : _GEN_6382; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6415 = 5'h4 == rd ? nzimm_C_LUI : _GEN_6383; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6416 = 5'h5 == rd ? nzimm_C_LUI : _GEN_6384; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6417 = 5'h6 == rd ? nzimm_C_LUI : _GEN_6385; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6418 = 5'h7 == rd ? nzimm_C_LUI : _GEN_6386; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6419 = 5'h8 == rd ? nzimm_C_LUI : _GEN_6387; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6420 = 5'h9 == rd ? nzimm_C_LUI : _GEN_6388; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6421 = 5'ha == rd ? nzimm_C_LUI : _GEN_6389; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6422 = 5'hb == rd ? nzimm_C_LUI : _GEN_6390; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6423 = 5'hc == rd ? nzimm_C_LUI : _GEN_6391; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6424 = 5'hd == rd ? nzimm_C_LUI : _GEN_6392; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6425 = 5'he == rd ? nzimm_C_LUI : _GEN_6393; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6426 = 5'hf == rd ? nzimm_C_LUI : _GEN_6394; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6427 = 5'h10 == rd ? nzimm_C_LUI : _GEN_6395; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6428 = 5'h11 == rd ? nzimm_C_LUI : _GEN_6396; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6429 = 5'h12 == rd ? nzimm_C_LUI : _GEN_6397; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6430 = 5'h13 == rd ? nzimm_C_LUI : _GEN_6398; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6431 = 5'h14 == rd ? nzimm_C_LUI : _GEN_6399; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6432 = 5'h15 == rd ? nzimm_C_LUI : _GEN_6400; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6433 = 5'h16 == rd ? nzimm_C_LUI : _GEN_6401; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6434 = 5'h17 == rd ? nzimm_C_LUI : _GEN_6402; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6435 = 5'h18 == rd ? nzimm_C_LUI : _GEN_6403; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6436 = 5'h19 == rd ? nzimm_C_LUI : _GEN_6404; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6437 = 5'h1a == rd ? nzimm_C_LUI : _GEN_6405; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6438 = 5'h1b == rd ? nzimm_C_LUI : _GEN_6406; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6439 = 5'h1c == rd ? nzimm_C_LUI : _GEN_6407; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6440 = 5'h1d == rd ? nzimm_C_LUI : _GEN_6408; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6441 = 5'h1e == rd ? nzimm_C_LUI : _GEN_6409; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6442 = 5'h1f == rd ? nzimm_C_LUI : _GEN_6410; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 212:{20,20}]
  wire [63:0] _GEN_6451 = _T_1146 ? _GEN_6412 : _GEN_6380; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6452 = _T_1146 ? _GEN_6413 : _GEN_6381; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6453 = _T_1146 ? _GEN_6414 : _GEN_6382; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6454 = _T_1146 ? _GEN_6415 : _GEN_6383; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6455 = _T_1146 ? _GEN_6416 : _GEN_6384; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6456 = _T_1146 ? _GEN_6417 : _GEN_6385; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6457 = _T_1146 ? _GEN_6418 : _GEN_6386; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6458 = _T_1146 ? _GEN_6419 : _GEN_6387; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6459 = _T_1146 ? _GEN_6420 : _GEN_6388; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6460 = _T_1146 ? _GEN_6421 : _GEN_6389; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6461 = _T_1146 ? _GEN_6422 : _GEN_6390; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6462 = _T_1146 ? _GEN_6423 : _GEN_6391; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6463 = _T_1146 ? _GEN_6424 : _GEN_6392; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6464 = _T_1146 ? _GEN_6425 : _GEN_6393; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6465 = _T_1146 ? _GEN_6426 : _GEN_6394; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6466 = _T_1146 ? _GEN_6427 : _GEN_6395; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6467 = _T_1146 ? _GEN_6428 : _GEN_6396; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6468 = _T_1146 ? _GEN_6429 : _GEN_6397; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6469 = _T_1146 ? _GEN_6430 : _GEN_6398; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6470 = _T_1146 ? _GEN_6431 : _GEN_6399; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6471 = _T_1146 ? _GEN_6432 : _GEN_6400; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6472 = _T_1146 ? _GEN_6433 : _GEN_6401; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6473 = _T_1146 ? _GEN_6434 : _GEN_6402; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6474 = _T_1146 ? _GEN_6435 : _GEN_6403; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6475 = _T_1146 ? _GEN_6436 : _GEN_6404; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6476 = _T_1146 ? _GEN_6437 : _GEN_6405; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6477 = _T_1146 ? _GEN_6438 : _GEN_6406; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6478 = _T_1146 ? _GEN_6439 : _GEN_6407; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6479 = _T_1146 ? _GEN_6440 : _GEN_6408; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6480 = _T_1146 ? _GEN_6441 : _GEN_6409; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6481 = _T_1146 ? _GEN_6442 : _GEN_6410; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 209:23]
  wire [63:0] _GEN_6483 = 5'h1 == rd ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6484 = 5'h2 == rd ? io_now_reg_2 : _GEN_6483; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6485 = 5'h3 == rd ? io_now_reg_3 : _GEN_6484; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6486 = 5'h4 == rd ? io_now_reg_4 : _GEN_6485; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6487 = 5'h5 == rd ? io_now_reg_5 : _GEN_6486; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6488 = 5'h6 == rd ? io_now_reg_6 : _GEN_6487; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6489 = 5'h7 == rd ? io_now_reg_7 : _GEN_6488; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6490 = 5'h8 == rd ? io_now_reg_8 : _GEN_6489; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6491 = 5'h9 == rd ? io_now_reg_9 : _GEN_6490; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6492 = 5'ha == rd ? io_now_reg_10 : _GEN_6491; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6493 = 5'hb == rd ? io_now_reg_11 : _GEN_6492; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6494 = 5'hc == rd ? io_now_reg_12 : _GEN_6493; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6495 = 5'hd == rd ? io_now_reg_13 : _GEN_6494; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6496 = 5'he == rd ? io_now_reg_14 : _GEN_6495; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6497 = 5'hf == rd ? io_now_reg_15 : _GEN_6496; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6498 = 5'h10 == rd ? io_now_reg_16 : _GEN_6497; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6499 = 5'h11 == rd ? io_now_reg_17 : _GEN_6498; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6500 = 5'h12 == rd ? io_now_reg_18 : _GEN_6499; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6501 = 5'h13 == rd ? io_now_reg_19 : _GEN_6500; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6502 = 5'h14 == rd ? io_now_reg_20 : _GEN_6501; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6503 = 5'h15 == rd ? io_now_reg_21 : _GEN_6502; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6504 = 5'h16 == rd ? io_now_reg_22 : _GEN_6503; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6505 = 5'h17 == rd ? io_now_reg_23 : _GEN_6504; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6506 = 5'h18 == rd ? io_now_reg_24 : _GEN_6505; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6507 = 5'h19 == rd ? io_now_reg_25 : _GEN_6506; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6508 = 5'h1a == rd ? io_now_reg_26 : _GEN_6507; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6509 = 5'h1b == rd ? io_now_reg_27 : _GEN_6508; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6510 = 5'h1c == rd ? io_now_reg_28 : _GEN_6509; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6511 = 5'h1d == rd ? io_now_reg_29 : _GEN_6510; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6512 = 5'h1e == rd ? io_now_reg_30 : _GEN_6511; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _GEN_6513 = 5'h1f == rd ? io_now_reg_31 : _GEN_6512; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{35,35}]
  wire [63:0] _next_reg_T_661 = _GEN_6513 + _imm_T_309; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:35]
  wire [63:0] _GEN_6515 = 5'h1 == rd ? _next_reg_T_661 : _GEN_6451; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6516 = 5'h2 == rd ? _next_reg_T_661 : _GEN_6452; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6517 = 5'h3 == rd ? _next_reg_T_661 : _GEN_6453; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6518 = 5'h4 == rd ? _next_reg_T_661 : _GEN_6454; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6519 = 5'h5 == rd ? _next_reg_T_661 : _GEN_6455; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6520 = 5'h6 == rd ? _next_reg_T_661 : _GEN_6456; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6521 = 5'h7 == rd ? _next_reg_T_661 : _GEN_6457; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6522 = 5'h8 == rd ? _next_reg_T_661 : _GEN_6458; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6523 = 5'h9 == rd ? _next_reg_T_661 : _GEN_6459; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6524 = 5'ha == rd ? _next_reg_T_661 : _GEN_6460; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6525 = 5'hb == rd ? _next_reg_T_661 : _GEN_6461; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6526 = 5'hc == rd ? _next_reg_T_661 : _GEN_6462; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6527 = 5'hd == rd ? _next_reg_T_661 : _GEN_6463; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6528 = 5'he == rd ? _next_reg_T_661 : _GEN_6464; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6529 = 5'hf == rd ? _next_reg_T_661 : _GEN_6465; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6530 = 5'h10 == rd ? _next_reg_T_661 : _GEN_6466; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6531 = 5'h11 == rd ? _next_reg_T_661 : _GEN_6467; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6532 = 5'h12 == rd ? _next_reg_T_661 : _GEN_6468; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6533 = 5'h13 == rd ? _next_reg_T_661 : _GEN_6469; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6534 = 5'h14 == rd ? _next_reg_T_661 : _GEN_6470; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6535 = 5'h15 == rd ? _next_reg_T_661 : _GEN_6471; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6536 = 5'h16 == rd ? _next_reg_T_661 : _GEN_6472; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6537 = 5'h17 == rd ? _next_reg_T_661 : _GEN_6473; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6538 = 5'h18 == rd ? _next_reg_T_661 : _GEN_6474; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6539 = 5'h19 == rd ? _next_reg_T_661 : _GEN_6475; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6540 = 5'h1a == rd ? _next_reg_T_661 : _GEN_6476; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6541 = 5'h1b == rd ? _next_reg_T_661 : _GEN_6477; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6542 = 5'h1c == rd ? _next_reg_T_661 : _GEN_6478; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6543 = 5'h1d == rd ? _next_reg_T_661 : _GEN_6479; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6544 = 5'h1e == rd ? _next_reg_T_661 : _GEN_6480; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6545 = 5'h1f == rd ? _next_reg_T_661 : _GEN_6481; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 218:{20,20}]
  wire [63:0] _GEN_6554 = _T_1161 ? _GEN_6515 : _GEN_6451; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6555 = _T_1161 ? _GEN_6516 : _GEN_6452; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6556 = _T_1161 ? _GEN_6517 : _GEN_6453; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6557 = _T_1161 ? _GEN_6518 : _GEN_6454; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6558 = _T_1161 ? _GEN_6519 : _GEN_6455; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6559 = _T_1161 ? _GEN_6520 : _GEN_6456; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6560 = _T_1161 ? _GEN_6521 : _GEN_6457; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6561 = _T_1161 ? _GEN_6522 : _GEN_6458; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6562 = _T_1161 ? _GEN_6523 : _GEN_6459; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6563 = _T_1161 ? _GEN_6524 : _GEN_6460; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6564 = _T_1161 ? _GEN_6525 : _GEN_6461; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6565 = _T_1161 ? _GEN_6526 : _GEN_6462; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6566 = _T_1161 ? _GEN_6527 : _GEN_6463; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6567 = _T_1161 ? _GEN_6528 : _GEN_6464; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6568 = _T_1161 ? _GEN_6529 : _GEN_6465; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6569 = _T_1161 ? _GEN_6530 : _GEN_6466; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6570 = _T_1161 ? _GEN_6531 : _GEN_6467; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6571 = _T_1161 ? _GEN_6532 : _GEN_6468; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6572 = _T_1161 ? _GEN_6533 : _GEN_6469; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6573 = _T_1161 ? _GEN_6534 : _GEN_6470; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6574 = _T_1161 ? _GEN_6535 : _GEN_6471; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6575 = _T_1161 ? _GEN_6536 : _GEN_6472; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6576 = _T_1161 ? _GEN_6537 : _GEN_6473; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6577 = _T_1161 ? _GEN_6538 : _GEN_6474; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6578 = _T_1161 ? _GEN_6539 : _GEN_6475; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6579 = _T_1161 ? _GEN_6540 : _GEN_6476; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6580 = _T_1161 ? _GEN_6541 : _GEN_6477; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6581 = _T_1161 ? _GEN_6542 : _GEN_6478; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6582 = _T_1161 ? _GEN_6543 : _GEN_6479; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6583 = _T_1161 ? _GEN_6544 : _GEN_6480; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [63:0] _GEN_6584 = _T_1161 ? _GEN_6545 : _GEN_6481; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 215:24]
  wire [9:0] _nzimm_C_ADDI16SP_T_7 = {inst[12],inst[4],inst[3],inst[5],inst[2],inst[6],4'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 85:10]
  wire  nzimm_C_ADDI16SP_signBit = _nzimm_C_ADDI16SP_T_7[9]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [53:0] _nzimm_C_ADDI16SP_T_9 = nzimm_C_ADDI16SP_signBit ? 54'h3fffffffffffff : 54'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] nzimm_C_ADDI16SP = {_nzimm_C_ADDI16SP_T_9,inst[12],inst[4],inst[3],inst[5],inst[2],inst[6],4'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _next_reg_2_T_1 = io_now_reg_2 + nzimm_C_ADDI16SP; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 223:37]
  wire [63:0] _GEN_6592 = _T_1173 ? _next_reg_2_T_1 : _GEN_6555; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 220:28 223:21]
  wire [63:0] nzimm_C_ADDI4SPN = {54'h0,inst[10],inst[9],inst[8],inst[7],inst[12],inst[11],inst[5],inst[6],2'h0}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [63:0] _next_reg_T_663 = io_now_reg_2 + nzimm_C_ADDI4SPN; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:44]
  wire [63:0] _GEN_6594 = 5'h1 == _T_1012 ? _next_reg_T_663 : _GEN_6554; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6595 = 5'h2 == _T_1012 ? _next_reg_T_663 : _GEN_6592; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6596 = 5'h3 == _T_1012 ? _next_reg_T_663 : _GEN_6556; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6597 = 5'h4 == _T_1012 ? _next_reg_T_663 : _GEN_6557; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6598 = 5'h5 == _T_1012 ? _next_reg_T_663 : _GEN_6558; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6599 = 5'h6 == _T_1012 ? _next_reg_T_663 : _GEN_6559; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6600 = 5'h7 == _T_1012 ? _next_reg_T_663 : _GEN_6560; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6601 = 5'h8 == _T_1012 ? _next_reg_T_663 : _GEN_6561; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6602 = 5'h9 == _T_1012 ? _next_reg_T_663 : _GEN_6562; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6603 = 5'ha == _T_1012 ? _next_reg_T_663 : _GEN_6563; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6604 = 5'hb == _T_1012 ? _next_reg_T_663 : _GEN_6564; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6605 = 5'hc == _T_1012 ? _next_reg_T_663 : _GEN_6565; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6606 = 5'hd == _T_1012 ? _next_reg_T_663 : _GEN_6566; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6607 = 5'he == _T_1012 ? _next_reg_T_663 : _GEN_6567; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6608 = 5'hf == _T_1012 ? _next_reg_T_663 : _GEN_6568; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6609 = 5'h10 == _T_1012 ? _next_reg_T_663 : _GEN_6569; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6610 = 5'h11 == _T_1012 ? _next_reg_T_663 : _GEN_6570; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6611 = 5'h12 == _T_1012 ? _next_reg_T_663 : _GEN_6571; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6612 = 5'h13 == _T_1012 ? _next_reg_T_663 : _GEN_6572; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6613 = 5'h14 == _T_1012 ? _next_reg_T_663 : _GEN_6573; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6614 = 5'h15 == _T_1012 ? _next_reg_T_663 : _GEN_6574; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6615 = 5'h16 == _T_1012 ? _next_reg_T_663 : _GEN_6575; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6616 = 5'h17 == _T_1012 ? _next_reg_T_663 : _GEN_6576; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6617 = 5'h18 == _T_1012 ? _next_reg_T_663 : _GEN_6577; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6618 = 5'h19 == _T_1012 ? _next_reg_T_663 : _GEN_6578; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6619 = 5'h1a == _T_1012 ? _next_reg_T_663 : _GEN_6579; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6620 = 5'h1b == _T_1012 ? _next_reg_T_663 : _GEN_6580; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6621 = 5'h1c == _T_1012 ? _next_reg_T_663 : _GEN_6581; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6622 = 5'h1d == _T_1012 ? _next_reg_T_663 : _GEN_6582; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6623 = 5'h1e == _T_1012 ? _next_reg_T_663 : _GEN_6583; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6624 = 5'h1f == _T_1012 ? _next_reg_T_663 : _GEN_6584; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 228:{28,28}]
  wire [63:0] _GEN_6631 = _T_1183 ? _GEN_6594 : _GEN_6554; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6632 = _T_1183 ? _GEN_6595 : _GEN_6592; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6633 = _T_1183 ? _GEN_6596 : _GEN_6556; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6634 = _T_1183 ? _GEN_6597 : _GEN_6557; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6635 = _T_1183 ? _GEN_6598 : _GEN_6558; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6636 = _T_1183 ? _GEN_6599 : _GEN_6559; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6637 = _T_1183 ? _GEN_6600 : _GEN_6560; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6638 = _T_1183 ? _GEN_6601 : _GEN_6561; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6639 = _T_1183 ? _GEN_6602 : _GEN_6562; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6640 = _T_1183 ? _GEN_6603 : _GEN_6563; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6641 = _T_1183 ? _GEN_6604 : _GEN_6564; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6642 = _T_1183 ? _GEN_6605 : _GEN_6565; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6643 = _T_1183 ? _GEN_6606 : _GEN_6566; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6644 = _T_1183 ? _GEN_6607 : _GEN_6567; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6645 = _T_1183 ? _GEN_6608 : _GEN_6568; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6646 = _T_1183 ? _GEN_6609 : _GEN_6569; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6647 = _T_1183 ? _GEN_6610 : _GEN_6570; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6648 = _T_1183 ? _GEN_6611 : _GEN_6571; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6649 = _T_1183 ? _GEN_6612 : _GEN_6572; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6650 = _T_1183 ? _GEN_6613 : _GEN_6573; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6651 = _T_1183 ? _GEN_6614 : _GEN_6574; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6652 = _T_1183 ? _GEN_6615 : _GEN_6575; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6653 = _T_1183 ? _GEN_6616 : _GEN_6576; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6654 = _T_1183 ? _GEN_6617 : _GEN_6577; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6655 = _T_1183 ? _GEN_6618 : _GEN_6578; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6656 = _T_1183 ? _GEN_6619 : _GEN_6579; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6657 = _T_1183 ? _GEN_6620 : _GEN_6580; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6658 = _T_1183 ? _GEN_6621 : _GEN_6581; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6659 = _T_1183 ? _GEN_6622 : _GEN_6582; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6660 = _T_1183 ? _GEN_6623 : _GEN_6583; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [63:0] _GEN_6661 = _T_1183 ? _GEN_6624 : _GEN_6584; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 225:28]
  wire [126:0] _GEN_6 = {{63'd0}, _GEN_6513}; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:35]
  wire [126:0] _next_reg_T_665 = _GEN_6 << imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:35]
  wire [63:0] _GEN_6663 = 5'h1 == rd ? _next_reg_T_665[63:0] : _GEN_6631; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6664 = 5'h2 == rd ? _next_reg_T_665[63:0] : _GEN_6632; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6665 = 5'h3 == rd ? _next_reg_T_665[63:0] : _GEN_6633; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6666 = 5'h4 == rd ? _next_reg_T_665[63:0] : _GEN_6634; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6667 = 5'h5 == rd ? _next_reg_T_665[63:0] : _GEN_6635; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6668 = 5'h6 == rd ? _next_reg_T_665[63:0] : _GEN_6636; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6669 = 5'h7 == rd ? _next_reg_T_665[63:0] : _GEN_6637; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6670 = 5'h8 == rd ? _next_reg_T_665[63:0] : _GEN_6638; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6671 = 5'h9 == rd ? _next_reg_T_665[63:0] : _GEN_6639; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6672 = 5'ha == rd ? _next_reg_T_665[63:0] : _GEN_6640; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6673 = 5'hb == rd ? _next_reg_T_665[63:0] : _GEN_6641; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6674 = 5'hc == rd ? _next_reg_T_665[63:0] : _GEN_6642; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6675 = 5'hd == rd ? _next_reg_T_665[63:0] : _GEN_6643; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6676 = 5'he == rd ? _next_reg_T_665[63:0] : _GEN_6644; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6677 = 5'hf == rd ? _next_reg_T_665[63:0] : _GEN_6645; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6678 = 5'h10 == rd ? _next_reg_T_665[63:0] : _GEN_6646; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6679 = 5'h11 == rd ? _next_reg_T_665[63:0] : _GEN_6647; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6680 = 5'h12 == rd ? _next_reg_T_665[63:0] : _GEN_6648; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6681 = 5'h13 == rd ? _next_reg_T_665[63:0] : _GEN_6649; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6682 = 5'h14 == rd ? _next_reg_T_665[63:0] : _GEN_6650; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6683 = 5'h15 == rd ? _next_reg_T_665[63:0] : _GEN_6651; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6684 = 5'h16 == rd ? _next_reg_T_665[63:0] : _GEN_6652; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6685 = 5'h17 == rd ? _next_reg_T_665[63:0] : _GEN_6653; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6686 = 5'h18 == rd ? _next_reg_T_665[63:0] : _GEN_6654; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6687 = 5'h19 == rd ? _next_reg_T_665[63:0] : _GEN_6655; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6688 = 5'h1a == rd ? _next_reg_T_665[63:0] : _GEN_6656; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6689 = 5'h1b == rd ? _next_reg_T_665[63:0] : _GEN_6657; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6690 = 5'h1c == rd ? _next_reg_T_665[63:0] : _GEN_6658; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6691 = 5'h1d == rd ? _next_reg_T_665[63:0] : _GEN_6659; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6692 = 5'h1e == rd ? _next_reg_T_665[63:0] : _GEN_6660; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6693 = 5'h1f == rd ? _next_reg_T_665[63:0] : _GEN_6661; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 233:{20,20}]
  wire [63:0] _GEN_6703 = _T_1199 ? _GEN_6663 : _GEN_6631; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6704 = _T_1199 ? _GEN_6664 : _GEN_6632; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6705 = _T_1199 ? _GEN_6665 : _GEN_6633; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6706 = _T_1199 ? _GEN_6666 : _GEN_6634; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6707 = _T_1199 ? _GEN_6667 : _GEN_6635; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6708 = _T_1199 ? _GEN_6668 : _GEN_6636; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6709 = _T_1199 ? _GEN_6669 : _GEN_6637; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6710 = _T_1199 ? _GEN_6670 : _GEN_6638; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6711 = _T_1199 ? _GEN_6671 : _GEN_6639; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6712 = _T_1199 ? _GEN_6672 : _GEN_6640; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6713 = _T_1199 ? _GEN_6673 : _GEN_6641; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6714 = _T_1199 ? _GEN_6674 : _GEN_6642; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6715 = _T_1199 ? _GEN_6675 : _GEN_6643; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6716 = _T_1199 ? _GEN_6676 : _GEN_6644; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6717 = _T_1199 ? _GEN_6677 : _GEN_6645; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6718 = _T_1199 ? _GEN_6678 : _GEN_6646; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6719 = _T_1199 ? _GEN_6679 : _GEN_6647; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6720 = _T_1199 ? _GEN_6680 : _GEN_6648; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6721 = _T_1199 ? _GEN_6681 : _GEN_6649; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6722 = _T_1199 ? _GEN_6682 : _GEN_6650; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6723 = _T_1199 ? _GEN_6683 : _GEN_6651; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6724 = _T_1199 ? _GEN_6684 : _GEN_6652; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6725 = _T_1199 ? _GEN_6685 : _GEN_6653; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6726 = _T_1199 ? _GEN_6686 : _GEN_6654; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6727 = _T_1199 ? _GEN_6687 : _GEN_6655; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6728 = _T_1199 ? _GEN_6688 : _GEN_6656; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6729 = _T_1199 ? _GEN_6689 : _GEN_6657; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6730 = _T_1199 ? _GEN_6690 : _GEN_6658; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6731 = _T_1199 ? _GEN_6691 : _GEN_6659; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6732 = _T_1199 ? _GEN_6692 : _GEN_6660; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6733 = _T_1199 ? _GEN_6693 : _GEN_6661; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 230:24]
  wire [63:0] _GEN_6735 = 5'h1 == _T_1012 ? io_now_reg_1 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6736 = 5'h2 == _T_1012 ? io_now_reg_2 : _GEN_6735; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6737 = 5'h3 == _T_1012 ? io_now_reg_3 : _GEN_6736; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6738 = 5'h4 == _T_1012 ? io_now_reg_4 : _GEN_6737; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6739 = 5'h5 == _T_1012 ? io_now_reg_5 : _GEN_6738; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6740 = 5'h6 == _T_1012 ? io_now_reg_6 : _GEN_6739; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6741 = 5'h7 == _T_1012 ? io_now_reg_7 : _GEN_6740; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6742 = 5'h8 == _T_1012 ? io_now_reg_8 : _GEN_6741; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6743 = 5'h9 == _T_1012 ? io_now_reg_9 : _GEN_6742; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6744 = 5'ha == _T_1012 ? io_now_reg_10 : _GEN_6743; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6745 = 5'hb == _T_1012 ? io_now_reg_11 : _GEN_6744; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6746 = 5'hc == _T_1012 ? io_now_reg_12 : _GEN_6745; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6747 = 5'hd == _T_1012 ? io_now_reg_13 : _GEN_6746; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6748 = 5'he == _T_1012 ? io_now_reg_14 : _GEN_6747; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6749 = 5'hf == _T_1012 ? io_now_reg_15 : _GEN_6748; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6750 = 5'h10 == _T_1012 ? io_now_reg_16 : _GEN_6749; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6751 = 5'h11 == _T_1012 ? io_now_reg_17 : _GEN_6750; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6752 = 5'h12 == _T_1012 ? io_now_reg_18 : _GEN_6751; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6753 = 5'h13 == _T_1012 ? io_now_reg_19 : _GEN_6752; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6754 = 5'h14 == _T_1012 ? io_now_reg_20 : _GEN_6753; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6755 = 5'h15 == _T_1012 ? io_now_reg_21 : _GEN_6754; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6756 = 5'h16 == _T_1012 ? io_now_reg_22 : _GEN_6755; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6757 = 5'h17 == _T_1012 ? io_now_reg_23 : _GEN_6756; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6758 = 5'h18 == _T_1012 ? io_now_reg_24 : _GEN_6757; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6759 = 5'h19 == _T_1012 ? io_now_reg_25 : _GEN_6758; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6760 = 5'h1a == _T_1012 ? io_now_reg_26 : _GEN_6759; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6761 = 5'h1b == _T_1012 ? io_now_reg_27 : _GEN_6760; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6762 = 5'h1c == _T_1012 ? io_now_reg_28 : _GEN_6761; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6763 = 5'h1d == _T_1012 ? io_now_reg_29 : _GEN_6762; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6764 = 5'h1e == _T_1012 ? io_now_reg_30 : _GEN_6763; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _GEN_6765 = 5'h1f == _T_1012 ? io_now_reg_31 : _GEN_6764; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{51,51}]
  wire [63:0] _next_reg_T_668 = _GEN_6765 >> imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:51]
  wire [63:0] _GEN_6767 = 5'h1 == _T_1012 ? _next_reg_T_668 : _GEN_6703; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6768 = 5'h2 == _T_1012 ? _next_reg_T_668 : _GEN_6704; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6769 = 5'h3 == _T_1012 ? _next_reg_T_668 : _GEN_6705; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6770 = 5'h4 == _T_1012 ? _next_reg_T_668 : _GEN_6706; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6771 = 5'h5 == _T_1012 ? _next_reg_T_668 : _GEN_6707; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6772 = 5'h6 == _T_1012 ? _next_reg_T_668 : _GEN_6708; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6773 = 5'h7 == _T_1012 ? _next_reg_T_668 : _GEN_6709; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6774 = 5'h8 == _T_1012 ? _next_reg_T_668 : _GEN_6710; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6775 = 5'h9 == _T_1012 ? _next_reg_T_668 : _GEN_6711; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6776 = 5'ha == _T_1012 ? _next_reg_T_668 : _GEN_6712; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6777 = 5'hb == _T_1012 ? _next_reg_T_668 : _GEN_6713; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6778 = 5'hc == _T_1012 ? _next_reg_T_668 : _GEN_6714; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6779 = 5'hd == _T_1012 ? _next_reg_T_668 : _GEN_6715; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6780 = 5'he == _T_1012 ? _next_reg_T_668 : _GEN_6716; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6781 = 5'hf == _T_1012 ? _next_reg_T_668 : _GEN_6717; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6782 = 5'h10 == _T_1012 ? _next_reg_T_668 : _GEN_6718; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6783 = 5'h11 == _T_1012 ? _next_reg_T_668 : _GEN_6719; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6784 = 5'h12 == _T_1012 ? _next_reg_T_668 : _GEN_6720; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6785 = 5'h13 == _T_1012 ? _next_reg_T_668 : _GEN_6721; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6786 = 5'h14 == _T_1012 ? _next_reg_T_668 : _GEN_6722; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6787 = 5'h15 == _T_1012 ? _next_reg_T_668 : _GEN_6723; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6788 = 5'h16 == _T_1012 ? _next_reg_T_668 : _GEN_6724; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6789 = 5'h17 == _T_1012 ? _next_reg_T_668 : _GEN_6725; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6790 = 5'h18 == _T_1012 ? _next_reg_T_668 : _GEN_6726; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6791 = 5'h19 == _T_1012 ? _next_reg_T_668 : _GEN_6727; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6792 = 5'h1a == _T_1012 ? _next_reg_T_668 : _GEN_6728; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6793 = 5'h1b == _T_1012 ? _next_reg_T_668 : _GEN_6729; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6794 = 5'h1c == _T_1012 ? _next_reg_T_668 : _GEN_6730; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6795 = 5'h1d == _T_1012 ? _next_reg_T_668 : _GEN_6731; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6796 = 5'h1e == _T_1012 ? _next_reg_T_668 : _GEN_6732; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6797 = 5'h1f == _T_1012 ? _next_reg_T_668 : _GEN_6733; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 238:{28,28}]
  wire [63:0] _GEN_6807 = _T_1212 ? _GEN_6767 : _GEN_6703; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6808 = _T_1212 ? _GEN_6768 : _GEN_6704; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6809 = _T_1212 ? _GEN_6769 : _GEN_6705; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6810 = _T_1212 ? _GEN_6770 : _GEN_6706; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6811 = _T_1212 ? _GEN_6771 : _GEN_6707; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6812 = _T_1212 ? _GEN_6772 : _GEN_6708; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6813 = _T_1212 ? _GEN_6773 : _GEN_6709; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6814 = _T_1212 ? _GEN_6774 : _GEN_6710; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6815 = _T_1212 ? _GEN_6775 : _GEN_6711; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6816 = _T_1212 ? _GEN_6776 : _GEN_6712; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6817 = _T_1212 ? _GEN_6777 : _GEN_6713; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6818 = _T_1212 ? _GEN_6778 : _GEN_6714; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6819 = _T_1212 ? _GEN_6779 : _GEN_6715; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6820 = _T_1212 ? _GEN_6780 : _GEN_6716; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6821 = _T_1212 ? _GEN_6781 : _GEN_6717; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6822 = _T_1212 ? _GEN_6782 : _GEN_6718; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6823 = _T_1212 ? _GEN_6783 : _GEN_6719; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6824 = _T_1212 ? _GEN_6784 : _GEN_6720; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6825 = _T_1212 ? _GEN_6785 : _GEN_6721; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6826 = _T_1212 ? _GEN_6786 : _GEN_6722; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6827 = _T_1212 ? _GEN_6787 : _GEN_6723; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6828 = _T_1212 ? _GEN_6788 : _GEN_6724; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6829 = _T_1212 ? _GEN_6789 : _GEN_6725; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6830 = _T_1212 ? _GEN_6790 : _GEN_6726; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6831 = _T_1212 ? _GEN_6791 : _GEN_6727; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6832 = _T_1212 ? _GEN_6792 : _GEN_6728; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6833 = _T_1212 ? _GEN_6793 : _GEN_6729; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6834 = _T_1212 ? _GEN_6794 : _GEN_6730; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6835 = _T_1212 ? _GEN_6795 : _GEN_6731; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6836 = _T_1212 ? _GEN_6796 : _GEN_6732; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _GEN_6837 = _T_1212 ? _GEN_6797 : _GEN_6733; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 235:24]
  wire [63:0] _next_reg_T_670 = 5'h1f == _T_1012 ? io_now_reg_31 : _GEN_6764; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:52]
  wire [63:0] _next_reg_T_673 = $signed(_next_reg_T_670) >>> imm[5:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:73]
  wire [63:0] _GEN_6871 = 5'h1 == _T_1012 ? _next_reg_T_673 : _GEN_6807; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6872 = 5'h2 == _T_1012 ? _next_reg_T_673 : _GEN_6808; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6873 = 5'h3 == _T_1012 ? _next_reg_T_673 : _GEN_6809; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6874 = 5'h4 == _T_1012 ? _next_reg_T_673 : _GEN_6810; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6875 = 5'h5 == _T_1012 ? _next_reg_T_673 : _GEN_6811; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6876 = 5'h6 == _T_1012 ? _next_reg_T_673 : _GEN_6812; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6877 = 5'h7 == _T_1012 ? _next_reg_T_673 : _GEN_6813; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6878 = 5'h8 == _T_1012 ? _next_reg_T_673 : _GEN_6814; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6879 = 5'h9 == _T_1012 ? _next_reg_T_673 : _GEN_6815; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6880 = 5'ha == _T_1012 ? _next_reg_T_673 : _GEN_6816; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6881 = 5'hb == _T_1012 ? _next_reg_T_673 : _GEN_6817; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6882 = 5'hc == _T_1012 ? _next_reg_T_673 : _GEN_6818; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6883 = 5'hd == _T_1012 ? _next_reg_T_673 : _GEN_6819; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6884 = 5'he == _T_1012 ? _next_reg_T_673 : _GEN_6820; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6885 = 5'hf == _T_1012 ? _next_reg_T_673 : _GEN_6821; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6886 = 5'h10 == _T_1012 ? _next_reg_T_673 : _GEN_6822; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6887 = 5'h11 == _T_1012 ? _next_reg_T_673 : _GEN_6823; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6888 = 5'h12 == _T_1012 ? _next_reg_T_673 : _GEN_6824; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6889 = 5'h13 == _T_1012 ? _next_reg_T_673 : _GEN_6825; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6890 = 5'h14 == _T_1012 ? _next_reg_T_673 : _GEN_6826; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6891 = 5'h15 == _T_1012 ? _next_reg_T_673 : _GEN_6827; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6892 = 5'h16 == _T_1012 ? _next_reg_T_673 : _GEN_6828; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6893 = 5'h17 == _T_1012 ? _next_reg_T_673 : _GEN_6829; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6894 = 5'h18 == _T_1012 ? _next_reg_T_673 : _GEN_6830; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6895 = 5'h19 == _T_1012 ? _next_reg_T_673 : _GEN_6831; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6896 = 5'h1a == _T_1012 ? _next_reg_T_673 : _GEN_6832; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6897 = 5'h1b == _T_1012 ? _next_reg_T_673 : _GEN_6833; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6898 = 5'h1c == _T_1012 ? _next_reg_T_673 : _GEN_6834; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6899 = 5'h1d == _T_1012 ? _next_reg_T_673 : _GEN_6835; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6900 = 5'h1e == _T_1012 ? _next_reg_T_673 : _GEN_6836; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6901 = 5'h1f == _T_1012 ? _next_reg_T_673 : _GEN_6837; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 243:{28,28}]
  wire [63:0] _GEN_6911 = _T_1226 ? _GEN_6871 : _GEN_6807; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6912 = _T_1226 ? _GEN_6872 : _GEN_6808; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6913 = _T_1226 ? _GEN_6873 : _GEN_6809; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6914 = _T_1226 ? _GEN_6874 : _GEN_6810; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6915 = _T_1226 ? _GEN_6875 : _GEN_6811; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6916 = _T_1226 ? _GEN_6876 : _GEN_6812; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6917 = _T_1226 ? _GEN_6877 : _GEN_6813; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6918 = _T_1226 ? _GEN_6878 : _GEN_6814; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6919 = _T_1226 ? _GEN_6879 : _GEN_6815; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6920 = _T_1226 ? _GEN_6880 : _GEN_6816; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6921 = _T_1226 ? _GEN_6881 : _GEN_6817; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6922 = _T_1226 ? _GEN_6882 : _GEN_6818; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6923 = _T_1226 ? _GEN_6883 : _GEN_6819; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6924 = _T_1226 ? _GEN_6884 : _GEN_6820; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6925 = _T_1226 ? _GEN_6885 : _GEN_6821; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6926 = _T_1226 ? _GEN_6886 : _GEN_6822; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6927 = _T_1226 ? _GEN_6887 : _GEN_6823; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6928 = _T_1226 ? _GEN_6888 : _GEN_6824; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6929 = _T_1226 ? _GEN_6889 : _GEN_6825; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6930 = _T_1226 ? _GEN_6890 : _GEN_6826; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6931 = _T_1226 ? _GEN_6891 : _GEN_6827; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6932 = _T_1226 ? _GEN_6892 : _GEN_6828; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6933 = _T_1226 ? _GEN_6893 : _GEN_6829; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6934 = _T_1226 ? _GEN_6894 : _GEN_6830; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6935 = _T_1226 ? _GEN_6895 : _GEN_6831; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6936 = _T_1226 ? _GEN_6896 : _GEN_6832; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6937 = _T_1226 ? _GEN_6897 : _GEN_6833; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6938 = _T_1226 ? _GEN_6898 : _GEN_6834; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6939 = _T_1226 ? _GEN_6899 : _GEN_6835; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6940 = _T_1226 ? _GEN_6900 : _GEN_6836; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _GEN_6941 = _T_1226 ? _GEN_6901 : _GEN_6837; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 240:24]
  wire [63:0] _next_reg_T_675 = _GEN_6765 & imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:51]
  wire [63:0] _GEN_6975 = 5'h1 == _T_1012 ? _next_reg_T_675 : _GEN_6911; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6976 = 5'h2 == _T_1012 ? _next_reg_T_675 : _GEN_6912; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6977 = 5'h3 == _T_1012 ? _next_reg_T_675 : _GEN_6913; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6978 = 5'h4 == _T_1012 ? _next_reg_T_675 : _GEN_6914; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6979 = 5'h5 == _T_1012 ? _next_reg_T_675 : _GEN_6915; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6980 = 5'h6 == _T_1012 ? _next_reg_T_675 : _GEN_6916; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6981 = 5'h7 == _T_1012 ? _next_reg_T_675 : _GEN_6917; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6982 = 5'h8 == _T_1012 ? _next_reg_T_675 : _GEN_6918; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6983 = 5'h9 == _T_1012 ? _next_reg_T_675 : _GEN_6919; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6984 = 5'ha == _T_1012 ? _next_reg_T_675 : _GEN_6920; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6985 = 5'hb == _T_1012 ? _next_reg_T_675 : _GEN_6921; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6986 = 5'hc == _T_1012 ? _next_reg_T_675 : _GEN_6922; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6987 = 5'hd == _T_1012 ? _next_reg_T_675 : _GEN_6923; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6988 = 5'he == _T_1012 ? _next_reg_T_675 : _GEN_6924; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6989 = 5'hf == _T_1012 ? _next_reg_T_675 : _GEN_6925; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6990 = 5'h10 == _T_1012 ? _next_reg_T_675 : _GEN_6926; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6991 = 5'h11 == _T_1012 ? _next_reg_T_675 : _GEN_6927; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6992 = 5'h12 == _T_1012 ? _next_reg_T_675 : _GEN_6928; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6993 = 5'h13 == _T_1012 ? _next_reg_T_675 : _GEN_6929; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6994 = 5'h14 == _T_1012 ? _next_reg_T_675 : _GEN_6930; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6995 = 5'h15 == _T_1012 ? _next_reg_T_675 : _GEN_6931; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6996 = 5'h16 == _T_1012 ? _next_reg_T_675 : _GEN_6932; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6997 = 5'h17 == _T_1012 ? _next_reg_T_675 : _GEN_6933; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6998 = 5'h18 == _T_1012 ? _next_reg_T_675 : _GEN_6934; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_6999 = 5'h19 == _T_1012 ? _next_reg_T_675 : _GEN_6935; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_7000 = 5'h1a == _T_1012 ? _next_reg_T_675 : _GEN_6936; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_7001 = 5'h1b == _T_1012 ? _next_reg_T_675 : _GEN_6937; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_7002 = 5'h1c == _T_1012 ? _next_reg_T_675 : _GEN_6938; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_7003 = 5'h1d == _T_1012 ? _next_reg_T_675 : _GEN_6939; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_7004 = 5'h1e == _T_1012 ? _next_reg_T_675 : _GEN_6940; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_7005 = 5'h1f == _T_1012 ? _next_reg_T_675 : _GEN_6941; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 248:{28,28}]
  wire [63:0] _GEN_7015 = _T_1234 ? _GEN_6975 : _GEN_6911; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7016 = _T_1234 ? _GEN_6976 : _GEN_6912; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7017 = _T_1234 ? _GEN_6977 : _GEN_6913; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7018 = _T_1234 ? _GEN_6978 : _GEN_6914; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7019 = _T_1234 ? _GEN_6979 : _GEN_6915; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7020 = _T_1234 ? _GEN_6980 : _GEN_6916; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7021 = _T_1234 ? _GEN_6981 : _GEN_6917; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7022 = _T_1234 ? _GEN_6982 : _GEN_6918; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7023 = _T_1234 ? _GEN_6983 : _GEN_6919; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7024 = _T_1234 ? _GEN_6984 : _GEN_6920; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7025 = _T_1234 ? _GEN_6985 : _GEN_6921; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7026 = _T_1234 ? _GEN_6986 : _GEN_6922; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7027 = _T_1234 ? _GEN_6987 : _GEN_6923; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7028 = _T_1234 ? _GEN_6988 : _GEN_6924; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7029 = _T_1234 ? _GEN_6989 : _GEN_6925; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7030 = _T_1234 ? _GEN_6990 : _GEN_6926; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7031 = _T_1234 ? _GEN_6991 : _GEN_6927; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7032 = _T_1234 ? _GEN_6992 : _GEN_6928; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7033 = _T_1234 ? _GEN_6993 : _GEN_6929; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7034 = _T_1234 ? _GEN_6994 : _GEN_6930; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7035 = _T_1234 ? _GEN_6995 : _GEN_6931; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7036 = _T_1234 ? _GEN_6996 : _GEN_6932; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7037 = _T_1234 ? _GEN_6997 : _GEN_6933; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7038 = _T_1234 ? _GEN_6998 : _GEN_6934; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7039 = _T_1234 ? _GEN_6999 : _GEN_6935; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7040 = _T_1234 ? _GEN_7000 : _GEN_6936; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7041 = _T_1234 ? _GEN_7001 : _GEN_6937; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7042 = _T_1234 ? _GEN_7002 : _GEN_6938; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7043 = _T_1234 ? _GEN_7003 : _GEN_6939; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7044 = _T_1234 ? _GEN_7004 : _GEN_6940; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _GEN_7045 = _T_1234 ? _GEN_7005 : _GEN_6941; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 245:24]
  wire [63:0] _next_reg_T_677 = io_now_reg_0 + _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:64]
  wire [63:0] _GEN_7047 = 5'h1 == rd ? _next_reg_T_677 : _GEN_7015; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7048 = 5'h2 == rd ? _next_reg_T_677 : _GEN_7016; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7049 = 5'h3 == rd ? _next_reg_T_677 : _GEN_7017; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7050 = 5'h4 == rd ? _next_reg_T_677 : _GEN_7018; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7051 = 5'h5 == rd ? _next_reg_T_677 : _GEN_7019; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7052 = 5'h6 == rd ? _next_reg_T_677 : _GEN_7020; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7053 = 5'h7 == rd ? _next_reg_T_677 : _GEN_7021; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7054 = 5'h8 == rd ? _next_reg_T_677 : _GEN_7022; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7055 = 5'h9 == rd ? _next_reg_T_677 : _GEN_7023; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7056 = 5'ha == rd ? _next_reg_T_677 : _GEN_7024; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7057 = 5'hb == rd ? _next_reg_T_677 : _GEN_7025; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7058 = 5'hc == rd ? _next_reg_T_677 : _GEN_7026; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7059 = 5'hd == rd ? _next_reg_T_677 : _GEN_7027; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7060 = 5'he == rd ? _next_reg_T_677 : _GEN_7028; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7061 = 5'hf == rd ? _next_reg_T_677 : _GEN_7029; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7062 = 5'h10 == rd ? _next_reg_T_677 : _GEN_7030; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7063 = 5'h11 == rd ? _next_reg_T_677 : _GEN_7031; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7064 = 5'h12 == rd ? _next_reg_T_677 : _GEN_7032; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7065 = 5'h13 == rd ? _next_reg_T_677 : _GEN_7033; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7066 = 5'h14 == rd ? _next_reg_T_677 : _GEN_7034; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7067 = 5'h15 == rd ? _next_reg_T_677 : _GEN_7035; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7068 = 5'h16 == rd ? _next_reg_T_677 : _GEN_7036; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7069 = 5'h17 == rd ? _next_reg_T_677 : _GEN_7037; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7070 = 5'h18 == rd ? _next_reg_T_677 : _GEN_7038; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7071 = 5'h19 == rd ? _next_reg_T_677 : _GEN_7039; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7072 = 5'h1a == rd ? _next_reg_T_677 : _GEN_7040; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7073 = 5'h1b == rd ? _next_reg_T_677 : _GEN_7041; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7074 = 5'h1c == rd ? _next_reg_T_677 : _GEN_7042; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7075 = 5'h1d == rd ? _next_reg_T_677 : _GEN_7043; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7076 = 5'h1e == rd ? _next_reg_T_677 : _GEN_7044; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7077 = 5'h1f == rd ? _next_reg_T_677 : _GEN_7045; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:{48,48}]
  wire [63:0] _GEN_7085 = _T_1248 ? _GEN_7047 : _GEN_7015; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7086 = _T_1248 ? _GEN_7048 : _GEN_7016; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7087 = _T_1248 ? _GEN_7049 : _GEN_7017; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7088 = _T_1248 ? _GEN_7050 : _GEN_7018; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7089 = _T_1248 ? _GEN_7051 : _GEN_7019; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7090 = _T_1248 ? _GEN_7052 : _GEN_7020; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7091 = _T_1248 ? _GEN_7053 : _GEN_7021; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7092 = _T_1248 ? _GEN_7054 : _GEN_7022; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7093 = _T_1248 ? _GEN_7055 : _GEN_7023; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7094 = _T_1248 ? _GEN_7056 : _GEN_7024; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7095 = _T_1248 ? _GEN_7057 : _GEN_7025; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7096 = _T_1248 ? _GEN_7058 : _GEN_7026; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7097 = _T_1248 ? _GEN_7059 : _GEN_7027; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7098 = _T_1248 ? _GEN_7060 : _GEN_7028; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7099 = _T_1248 ? _GEN_7061 : _GEN_7029; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7100 = _T_1248 ? _GEN_7062 : _GEN_7030; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7101 = _T_1248 ? _GEN_7063 : _GEN_7031; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7102 = _T_1248 ? _GEN_7064 : _GEN_7032; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7103 = _T_1248 ? _GEN_7065 : _GEN_7033; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7104 = _T_1248 ? _GEN_7066 : _GEN_7034; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7105 = _T_1248 ? _GEN_7067 : _GEN_7035; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7106 = _T_1248 ? _GEN_7068 : _GEN_7036; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7107 = _T_1248 ? _GEN_7069 : _GEN_7037; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7108 = _T_1248 ? _GEN_7070 : _GEN_7038; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7109 = _T_1248 ? _GEN_7071 : _GEN_7039; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7110 = _T_1248 ? _GEN_7072 : _GEN_7040; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7111 = _T_1248 ? _GEN_7073 : _GEN_7041; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7112 = _T_1248 ? _GEN_7074 : _GEN_7042; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7113 = _T_1248 ? _GEN_7075 : _GEN_7043; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7114 = _T_1248 ? _GEN_7076 : _GEN_7044; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _GEN_7115 = _T_1248 ? _GEN_7077 : _GEN_7045; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 251:23]
  wire [63:0] _next_reg_T_679 = _GEN_6513 + _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:63]
  wire [63:0] _GEN_7117 = 5'h1 == rd ? _next_reg_T_679 : _GEN_7085; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7118 = 5'h2 == rd ? _next_reg_T_679 : _GEN_7086; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7119 = 5'h3 == rd ? _next_reg_T_679 : _GEN_7087; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7120 = 5'h4 == rd ? _next_reg_T_679 : _GEN_7088; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7121 = 5'h5 == rd ? _next_reg_T_679 : _GEN_7089; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7122 = 5'h6 == rd ? _next_reg_T_679 : _GEN_7090; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7123 = 5'h7 == rd ? _next_reg_T_679 : _GEN_7091; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7124 = 5'h8 == rd ? _next_reg_T_679 : _GEN_7092; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7125 = 5'h9 == rd ? _next_reg_T_679 : _GEN_7093; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7126 = 5'ha == rd ? _next_reg_T_679 : _GEN_7094; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7127 = 5'hb == rd ? _next_reg_T_679 : _GEN_7095; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7128 = 5'hc == rd ? _next_reg_T_679 : _GEN_7096; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7129 = 5'hd == rd ? _next_reg_T_679 : _GEN_7097; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7130 = 5'he == rd ? _next_reg_T_679 : _GEN_7098; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7131 = 5'hf == rd ? _next_reg_T_679 : _GEN_7099; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7132 = 5'h10 == rd ? _next_reg_T_679 : _GEN_7100; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7133 = 5'h11 == rd ? _next_reg_T_679 : _GEN_7101; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7134 = 5'h12 == rd ? _next_reg_T_679 : _GEN_7102; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7135 = 5'h13 == rd ? _next_reg_T_679 : _GEN_7103; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7136 = 5'h14 == rd ? _next_reg_T_679 : _GEN_7104; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7137 = 5'h15 == rd ? _next_reg_T_679 : _GEN_7105; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7138 = 5'h16 == rd ? _next_reg_T_679 : _GEN_7106; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7139 = 5'h17 == rd ? _next_reg_T_679 : _GEN_7107; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7140 = 5'h18 == rd ? _next_reg_T_679 : _GEN_7108; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7141 = 5'h19 == rd ? _next_reg_T_679 : _GEN_7109; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7142 = 5'h1a == rd ? _next_reg_T_679 : _GEN_7110; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7143 = 5'h1b == rd ? _next_reg_T_679 : _GEN_7111; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7144 = 5'h1c == rd ? _next_reg_T_679 : _GEN_7112; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7145 = 5'h1d == rd ? _next_reg_T_679 : _GEN_7113; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7146 = 5'h1e == rd ? _next_reg_T_679 : _GEN_7114; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7147 = 5'h1f == rd ? _next_reg_T_679 : _GEN_7115; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:{48,48}]
  wire [63:0] _GEN_7155 = _T_1260 ? _GEN_7117 : _GEN_7085; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7156 = _T_1260 ? _GEN_7118 : _GEN_7086; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7157 = _T_1260 ? _GEN_7119 : _GEN_7087; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7158 = _T_1260 ? _GEN_7120 : _GEN_7088; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7159 = _T_1260 ? _GEN_7121 : _GEN_7089; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7160 = _T_1260 ? _GEN_7122 : _GEN_7090; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7161 = _T_1260 ? _GEN_7123 : _GEN_7091; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7162 = _T_1260 ? _GEN_7124 : _GEN_7092; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7163 = _T_1260 ? _GEN_7125 : _GEN_7093; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7164 = _T_1260 ? _GEN_7126 : _GEN_7094; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7165 = _T_1260 ? _GEN_7127 : _GEN_7095; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7166 = _T_1260 ? _GEN_7128 : _GEN_7096; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7167 = _T_1260 ? _GEN_7129 : _GEN_7097; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7168 = _T_1260 ? _GEN_7130 : _GEN_7098; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7169 = _T_1260 ? _GEN_7131 : _GEN_7099; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7170 = _T_1260 ? _GEN_7132 : _GEN_7100; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7171 = _T_1260 ? _GEN_7133 : _GEN_7101; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7172 = _T_1260 ? _GEN_7134 : _GEN_7102; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7173 = _T_1260 ? _GEN_7135 : _GEN_7103; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7174 = _T_1260 ? _GEN_7136 : _GEN_7104; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7175 = _T_1260 ? _GEN_7137 : _GEN_7105; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7176 = _T_1260 ? _GEN_7138 : _GEN_7106; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7177 = _T_1260 ? _GEN_7139 : _GEN_7107; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7178 = _T_1260 ? _GEN_7140 : _GEN_7108; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7179 = _T_1260 ? _GEN_7141 : _GEN_7109; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7180 = _T_1260 ? _GEN_7142 : _GEN_7110; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7181 = _T_1260 ? _GEN_7143 : _GEN_7111; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7182 = _T_1260 ? _GEN_7144 : _GEN_7112; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7183 = _T_1260 ? _GEN_7145 : _GEN_7113; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7184 = _T_1260 ? _GEN_7146 : _GEN_7114; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _GEN_7185 = _T_1260 ? _GEN_7147 : _GEN_7115; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 252:23]
  wire [63:0] _next_reg_T_682 = _GEN_6765 & _GEN_6191; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:79]
  wire [63:0] _GEN_7251 = 5'h1 == _T_1012 ? _next_reg_T_682 : _GEN_7155; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7252 = 5'h2 == _T_1012 ? _next_reg_T_682 : _GEN_7156; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7253 = 5'h3 == _T_1012 ? _next_reg_T_682 : _GEN_7157; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7254 = 5'h4 == _T_1012 ? _next_reg_T_682 : _GEN_7158; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7255 = 5'h5 == _T_1012 ? _next_reg_T_682 : _GEN_7159; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7256 = 5'h6 == _T_1012 ? _next_reg_T_682 : _GEN_7160; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7257 = 5'h7 == _T_1012 ? _next_reg_T_682 : _GEN_7161; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7258 = 5'h8 == _T_1012 ? _next_reg_T_682 : _GEN_7162; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7259 = 5'h9 == _T_1012 ? _next_reg_T_682 : _GEN_7163; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7260 = 5'ha == _T_1012 ? _next_reg_T_682 : _GEN_7164; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7261 = 5'hb == _T_1012 ? _next_reg_T_682 : _GEN_7165; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7262 = 5'hc == _T_1012 ? _next_reg_T_682 : _GEN_7166; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7263 = 5'hd == _T_1012 ? _next_reg_T_682 : _GEN_7167; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7264 = 5'he == _T_1012 ? _next_reg_T_682 : _GEN_7168; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7265 = 5'hf == _T_1012 ? _next_reg_T_682 : _GEN_7169; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7266 = 5'h10 == _T_1012 ? _next_reg_T_682 : _GEN_7170; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7267 = 5'h11 == _T_1012 ? _next_reg_T_682 : _GEN_7171; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7268 = 5'h12 == _T_1012 ? _next_reg_T_682 : _GEN_7172; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7269 = 5'h13 == _T_1012 ? _next_reg_T_682 : _GEN_7173; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7270 = 5'h14 == _T_1012 ? _next_reg_T_682 : _GEN_7174; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7271 = 5'h15 == _T_1012 ? _next_reg_T_682 : _GEN_7175; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7272 = 5'h16 == _T_1012 ? _next_reg_T_682 : _GEN_7176; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7273 = 5'h17 == _T_1012 ? _next_reg_T_682 : _GEN_7177; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7274 = 5'h18 == _T_1012 ? _next_reg_T_682 : _GEN_7178; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7275 = 5'h19 == _T_1012 ? _next_reg_T_682 : _GEN_7179; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7276 = 5'h1a == _T_1012 ? _next_reg_T_682 : _GEN_7180; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7277 = 5'h1b == _T_1012 ? _next_reg_T_682 : _GEN_7181; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7278 = 5'h1c == _T_1012 ? _next_reg_T_682 : _GEN_7182; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7279 = 5'h1d == _T_1012 ? _next_reg_T_682 : _GEN_7183; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7280 = 5'h1e == _T_1012 ? _next_reg_T_682 : _GEN_7184; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7281 = 5'h1f == _T_1012 ? _next_reg_T_682 : _GEN_7185; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:{56,56}]
  wire [63:0] _GEN_7290 = _T_1266 ? _GEN_7251 : _GEN_7155; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7291 = _T_1266 ? _GEN_7252 : _GEN_7156; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7292 = _T_1266 ? _GEN_7253 : _GEN_7157; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7293 = _T_1266 ? _GEN_7254 : _GEN_7158; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7294 = _T_1266 ? _GEN_7255 : _GEN_7159; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7295 = _T_1266 ? _GEN_7256 : _GEN_7160; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7296 = _T_1266 ? _GEN_7257 : _GEN_7161; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7297 = _T_1266 ? _GEN_7258 : _GEN_7162; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7298 = _T_1266 ? _GEN_7259 : _GEN_7163; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7299 = _T_1266 ? _GEN_7260 : _GEN_7164; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7300 = _T_1266 ? _GEN_7261 : _GEN_7165; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7301 = _T_1266 ? _GEN_7262 : _GEN_7166; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7302 = _T_1266 ? _GEN_7263 : _GEN_7167; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7303 = _T_1266 ? _GEN_7264 : _GEN_7168; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7304 = _T_1266 ? _GEN_7265 : _GEN_7169; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7305 = _T_1266 ? _GEN_7266 : _GEN_7170; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7306 = _T_1266 ? _GEN_7267 : _GEN_7171; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7307 = _T_1266 ? _GEN_7268 : _GEN_7172; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7308 = _T_1266 ? _GEN_7269 : _GEN_7173; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7309 = _T_1266 ? _GEN_7270 : _GEN_7174; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7310 = _T_1266 ? _GEN_7271 : _GEN_7175; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7311 = _T_1266 ? _GEN_7272 : _GEN_7176; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7312 = _T_1266 ? _GEN_7273 : _GEN_7177; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7313 = _T_1266 ? _GEN_7274 : _GEN_7178; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7314 = _T_1266 ? _GEN_7275 : _GEN_7179; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7315 = _T_1266 ? _GEN_7276 : _GEN_7180; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7316 = _T_1266 ? _GEN_7277 : _GEN_7181; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7317 = _T_1266 ? _GEN_7278 : _GEN_7182; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7318 = _T_1266 ? _GEN_7279 : _GEN_7183; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7319 = _T_1266 ? _GEN_7280 : _GEN_7184; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _GEN_7320 = _T_1266 ? _GEN_7281 : _GEN_7185; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 253:23]
  wire [63:0] _next_reg_T_685 = _GEN_6765 | _GEN_6191; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:79]
  wire [63:0] _GEN_7386 = 5'h1 == _T_1012 ? _next_reg_T_685 : _GEN_7290; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7387 = 5'h2 == _T_1012 ? _next_reg_T_685 : _GEN_7291; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7388 = 5'h3 == _T_1012 ? _next_reg_T_685 : _GEN_7292; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7389 = 5'h4 == _T_1012 ? _next_reg_T_685 : _GEN_7293; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7390 = 5'h5 == _T_1012 ? _next_reg_T_685 : _GEN_7294; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7391 = 5'h6 == _T_1012 ? _next_reg_T_685 : _GEN_7295; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7392 = 5'h7 == _T_1012 ? _next_reg_T_685 : _GEN_7296; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7393 = 5'h8 == _T_1012 ? _next_reg_T_685 : _GEN_7297; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7394 = 5'h9 == _T_1012 ? _next_reg_T_685 : _GEN_7298; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7395 = 5'ha == _T_1012 ? _next_reg_T_685 : _GEN_7299; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7396 = 5'hb == _T_1012 ? _next_reg_T_685 : _GEN_7300; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7397 = 5'hc == _T_1012 ? _next_reg_T_685 : _GEN_7301; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7398 = 5'hd == _T_1012 ? _next_reg_T_685 : _GEN_7302; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7399 = 5'he == _T_1012 ? _next_reg_T_685 : _GEN_7303; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7400 = 5'hf == _T_1012 ? _next_reg_T_685 : _GEN_7304; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7401 = 5'h10 == _T_1012 ? _next_reg_T_685 : _GEN_7305; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7402 = 5'h11 == _T_1012 ? _next_reg_T_685 : _GEN_7306; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7403 = 5'h12 == _T_1012 ? _next_reg_T_685 : _GEN_7307; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7404 = 5'h13 == _T_1012 ? _next_reg_T_685 : _GEN_7308; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7405 = 5'h14 == _T_1012 ? _next_reg_T_685 : _GEN_7309; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7406 = 5'h15 == _T_1012 ? _next_reg_T_685 : _GEN_7310; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7407 = 5'h16 == _T_1012 ? _next_reg_T_685 : _GEN_7311; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7408 = 5'h17 == _T_1012 ? _next_reg_T_685 : _GEN_7312; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7409 = 5'h18 == _T_1012 ? _next_reg_T_685 : _GEN_7313; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7410 = 5'h19 == _T_1012 ? _next_reg_T_685 : _GEN_7314; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7411 = 5'h1a == _T_1012 ? _next_reg_T_685 : _GEN_7315; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7412 = 5'h1b == _T_1012 ? _next_reg_T_685 : _GEN_7316; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7413 = 5'h1c == _T_1012 ? _next_reg_T_685 : _GEN_7317; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7414 = 5'h1d == _T_1012 ? _next_reg_T_685 : _GEN_7318; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7415 = 5'h1e == _T_1012 ? _next_reg_T_685 : _GEN_7319; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7416 = 5'h1f == _T_1012 ? _next_reg_T_685 : _GEN_7320; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:{56,56}]
  wire [63:0] _GEN_7425 = _T_1274 ? _GEN_7386 : _GEN_7290; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7426 = _T_1274 ? _GEN_7387 : _GEN_7291; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7427 = _T_1274 ? _GEN_7388 : _GEN_7292; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7428 = _T_1274 ? _GEN_7389 : _GEN_7293; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7429 = _T_1274 ? _GEN_7390 : _GEN_7294; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7430 = _T_1274 ? _GEN_7391 : _GEN_7295; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7431 = _T_1274 ? _GEN_7392 : _GEN_7296; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7432 = _T_1274 ? _GEN_7393 : _GEN_7297; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7433 = _T_1274 ? _GEN_7394 : _GEN_7298; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7434 = _T_1274 ? _GEN_7395 : _GEN_7299; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7435 = _T_1274 ? _GEN_7396 : _GEN_7300; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7436 = _T_1274 ? _GEN_7397 : _GEN_7301; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7437 = _T_1274 ? _GEN_7398 : _GEN_7302; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7438 = _T_1274 ? _GEN_7399 : _GEN_7303; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7439 = _T_1274 ? _GEN_7400 : _GEN_7304; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7440 = _T_1274 ? _GEN_7401 : _GEN_7305; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7441 = _T_1274 ? _GEN_7402 : _GEN_7306; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7442 = _T_1274 ? _GEN_7403 : _GEN_7307; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7443 = _T_1274 ? _GEN_7404 : _GEN_7308; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7444 = _T_1274 ? _GEN_7405 : _GEN_7309; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7445 = _T_1274 ? _GEN_7406 : _GEN_7310; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7446 = _T_1274 ? _GEN_7407 : _GEN_7311; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7447 = _T_1274 ? _GEN_7408 : _GEN_7312; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7448 = _T_1274 ? _GEN_7409 : _GEN_7313; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7449 = _T_1274 ? _GEN_7410 : _GEN_7314; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7450 = _T_1274 ? _GEN_7411 : _GEN_7315; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7451 = _T_1274 ? _GEN_7412 : _GEN_7316; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7452 = _T_1274 ? _GEN_7413 : _GEN_7317; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7453 = _T_1274 ? _GEN_7414 : _GEN_7318; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7454 = _T_1274 ? _GEN_7415 : _GEN_7319; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _GEN_7455 = _T_1274 ? _GEN_7416 : _GEN_7320; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 254:23]
  wire [63:0] _next_reg_T_688 = _GEN_6765 ^ _GEN_6191; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:79]
  wire [63:0] _GEN_7521 = 5'h1 == _T_1012 ? _next_reg_T_688 : _GEN_7425; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7522 = 5'h2 == _T_1012 ? _next_reg_T_688 : _GEN_7426; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7523 = 5'h3 == _T_1012 ? _next_reg_T_688 : _GEN_7427; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7524 = 5'h4 == _T_1012 ? _next_reg_T_688 : _GEN_7428; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7525 = 5'h5 == _T_1012 ? _next_reg_T_688 : _GEN_7429; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7526 = 5'h6 == _T_1012 ? _next_reg_T_688 : _GEN_7430; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7527 = 5'h7 == _T_1012 ? _next_reg_T_688 : _GEN_7431; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7528 = 5'h8 == _T_1012 ? _next_reg_T_688 : _GEN_7432; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7529 = 5'h9 == _T_1012 ? _next_reg_T_688 : _GEN_7433; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7530 = 5'ha == _T_1012 ? _next_reg_T_688 : _GEN_7434; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7531 = 5'hb == _T_1012 ? _next_reg_T_688 : _GEN_7435; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7532 = 5'hc == _T_1012 ? _next_reg_T_688 : _GEN_7436; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7533 = 5'hd == _T_1012 ? _next_reg_T_688 : _GEN_7437; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7534 = 5'he == _T_1012 ? _next_reg_T_688 : _GEN_7438; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7535 = 5'hf == _T_1012 ? _next_reg_T_688 : _GEN_7439; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7536 = 5'h10 == _T_1012 ? _next_reg_T_688 : _GEN_7440; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7537 = 5'h11 == _T_1012 ? _next_reg_T_688 : _GEN_7441; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7538 = 5'h12 == _T_1012 ? _next_reg_T_688 : _GEN_7442; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7539 = 5'h13 == _T_1012 ? _next_reg_T_688 : _GEN_7443; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7540 = 5'h14 == _T_1012 ? _next_reg_T_688 : _GEN_7444; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7541 = 5'h15 == _T_1012 ? _next_reg_T_688 : _GEN_7445; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7542 = 5'h16 == _T_1012 ? _next_reg_T_688 : _GEN_7446; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7543 = 5'h17 == _T_1012 ? _next_reg_T_688 : _GEN_7447; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7544 = 5'h18 == _T_1012 ? _next_reg_T_688 : _GEN_7448; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7545 = 5'h19 == _T_1012 ? _next_reg_T_688 : _GEN_7449; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7546 = 5'h1a == _T_1012 ? _next_reg_T_688 : _GEN_7450; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7547 = 5'h1b == _T_1012 ? _next_reg_T_688 : _GEN_7451; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7548 = 5'h1c == _T_1012 ? _next_reg_T_688 : _GEN_7452; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7549 = 5'h1d == _T_1012 ? _next_reg_T_688 : _GEN_7453; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7550 = 5'h1e == _T_1012 ? _next_reg_T_688 : _GEN_7454; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7551 = 5'h1f == _T_1012 ? _next_reg_T_688 : _GEN_7455; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:{56,56}]
  wire [63:0] _GEN_7560 = _T_1282 ? _GEN_7521 : _GEN_7425; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7561 = _T_1282 ? _GEN_7522 : _GEN_7426; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7562 = _T_1282 ? _GEN_7523 : _GEN_7427; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7563 = _T_1282 ? _GEN_7524 : _GEN_7428; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7564 = _T_1282 ? _GEN_7525 : _GEN_7429; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7565 = _T_1282 ? _GEN_7526 : _GEN_7430; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7566 = _T_1282 ? _GEN_7527 : _GEN_7431; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7567 = _T_1282 ? _GEN_7528 : _GEN_7432; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7568 = _T_1282 ? _GEN_7529 : _GEN_7433; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7569 = _T_1282 ? _GEN_7530 : _GEN_7434; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7570 = _T_1282 ? _GEN_7531 : _GEN_7435; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7571 = _T_1282 ? _GEN_7532 : _GEN_7436; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7572 = _T_1282 ? _GEN_7533 : _GEN_7437; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7573 = _T_1282 ? _GEN_7534 : _GEN_7438; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7574 = _T_1282 ? _GEN_7535 : _GEN_7439; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7575 = _T_1282 ? _GEN_7536 : _GEN_7440; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7576 = _T_1282 ? _GEN_7537 : _GEN_7441; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7577 = _T_1282 ? _GEN_7538 : _GEN_7442; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7578 = _T_1282 ? _GEN_7539 : _GEN_7443; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7579 = _T_1282 ? _GEN_7540 : _GEN_7444; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7580 = _T_1282 ? _GEN_7541 : _GEN_7445; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7581 = _T_1282 ? _GEN_7542 : _GEN_7446; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7582 = _T_1282 ? _GEN_7543 : _GEN_7447; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7583 = _T_1282 ? _GEN_7544 : _GEN_7448; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7584 = _T_1282 ? _GEN_7545 : _GEN_7449; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7585 = _T_1282 ? _GEN_7546 : _GEN_7450; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7586 = _T_1282 ? _GEN_7547 : _GEN_7451; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7587 = _T_1282 ? _GEN_7548 : _GEN_7452; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7588 = _T_1282 ? _GEN_7549 : _GEN_7453; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7589 = _T_1282 ? _GEN_7550 : _GEN_7454; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _GEN_7590 = _T_1282 ? _GEN_7551 : _GEN_7455; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 255:23]
  wire [63:0] _next_reg_T_692 = _GEN_6765 - _GEN_6191; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:79]
  wire [63:0] _GEN_7656 = 5'h1 == _T_1012 ? _next_reg_T_692 : _GEN_7560; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7657 = 5'h2 == _T_1012 ? _next_reg_T_692 : _GEN_7561; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7658 = 5'h3 == _T_1012 ? _next_reg_T_692 : _GEN_7562; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7659 = 5'h4 == _T_1012 ? _next_reg_T_692 : _GEN_7563; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7660 = 5'h5 == _T_1012 ? _next_reg_T_692 : _GEN_7564; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7661 = 5'h6 == _T_1012 ? _next_reg_T_692 : _GEN_7565; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7662 = 5'h7 == _T_1012 ? _next_reg_T_692 : _GEN_7566; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7663 = 5'h8 == _T_1012 ? _next_reg_T_692 : _GEN_7567; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7664 = 5'h9 == _T_1012 ? _next_reg_T_692 : _GEN_7568; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7665 = 5'ha == _T_1012 ? _next_reg_T_692 : _GEN_7569; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7666 = 5'hb == _T_1012 ? _next_reg_T_692 : _GEN_7570; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7667 = 5'hc == _T_1012 ? _next_reg_T_692 : _GEN_7571; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7668 = 5'hd == _T_1012 ? _next_reg_T_692 : _GEN_7572; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7669 = 5'he == _T_1012 ? _next_reg_T_692 : _GEN_7573; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7670 = 5'hf == _T_1012 ? _next_reg_T_692 : _GEN_7574; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7671 = 5'h10 == _T_1012 ? _next_reg_T_692 : _GEN_7575; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7672 = 5'h11 == _T_1012 ? _next_reg_T_692 : _GEN_7576; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7673 = 5'h12 == _T_1012 ? _next_reg_T_692 : _GEN_7577; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7674 = 5'h13 == _T_1012 ? _next_reg_T_692 : _GEN_7578; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7675 = 5'h14 == _T_1012 ? _next_reg_T_692 : _GEN_7579; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7676 = 5'h15 == _T_1012 ? _next_reg_T_692 : _GEN_7580; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7677 = 5'h16 == _T_1012 ? _next_reg_T_692 : _GEN_7581; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7678 = 5'h17 == _T_1012 ? _next_reg_T_692 : _GEN_7582; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7679 = 5'h18 == _T_1012 ? _next_reg_T_692 : _GEN_7583; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7680 = 5'h19 == _T_1012 ? _next_reg_T_692 : _GEN_7584; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7681 = 5'h1a == _T_1012 ? _next_reg_T_692 : _GEN_7585; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7682 = 5'h1b == _T_1012 ? _next_reg_T_692 : _GEN_7586; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7683 = 5'h1c == _T_1012 ? _next_reg_T_692 : _GEN_7587; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7684 = 5'h1d == _T_1012 ? _next_reg_T_692 : _GEN_7588; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7685 = 5'h1e == _T_1012 ? _next_reg_T_692 : _GEN_7589; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7686 = 5'h1f == _T_1012 ? _next_reg_T_692 : _GEN_7590; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:{56,56}]
  wire [63:0] _GEN_7695 = _T_1290 ? _GEN_7656 : _GEN_7560; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7696 = _T_1290 ? _GEN_7657 : _GEN_7561; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7697 = _T_1290 ? _GEN_7658 : _GEN_7562; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7698 = _T_1290 ? _GEN_7659 : _GEN_7563; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7699 = _T_1290 ? _GEN_7660 : _GEN_7564; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7700 = _T_1290 ? _GEN_7661 : _GEN_7565; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7701 = _T_1290 ? _GEN_7662 : _GEN_7566; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7702 = _T_1290 ? _GEN_7663 : _GEN_7567; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7703 = _T_1290 ? _GEN_7664 : _GEN_7568; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7704 = _T_1290 ? _GEN_7665 : _GEN_7569; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7705 = _T_1290 ? _GEN_7666 : _GEN_7570; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7706 = _T_1290 ? _GEN_7667 : _GEN_7571; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7707 = _T_1290 ? _GEN_7668 : _GEN_7572; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7708 = _T_1290 ? _GEN_7669 : _GEN_7573; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7709 = _T_1290 ? _GEN_7670 : _GEN_7574; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7710 = _T_1290 ? _GEN_7671 : _GEN_7575; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7711 = _T_1290 ? _GEN_7672 : _GEN_7576; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7712 = _T_1290 ? _GEN_7673 : _GEN_7577; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7713 = _T_1290 ? _GEN_7674 : _GEN_7578; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7714 = _T_1290 ? _GEN_7675 : _GEN_7579; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7715 = _T_1290 ? _GEN_7676 : _GEN_7580; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7716 = _T_1290 ? _GEN_7677 : _GEN_7581; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7717 = _T_1290 ? _GEN_7678 : _GEN_7582; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7718 = _T_1290 ? _GEN_7679 : _GEN_7583; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7719 = _T_1290 ? _GEN_7680 : _GEN_7584; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7720 = _T_1290 ? _GEN_7681 : _GEN_7585; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7721 = _T_1290 ? _GEN_7682 : _GEN_7586; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7722 = _T_1290 ? _GEN_7683 : _GEN_7587; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7723 = _T_1290 ? _GEN_7684 : _GEN_7588; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7724 = _T_1290 ? _GEN_7685 : _GEN_7589; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire [63:0] _GEN_7725 = _T_1290 ? _GEN_7686 : _GEN_7590; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 256:23]
  wire  _GEN_7756 = next_reg_LevelVec_10_1_valid | _GEN_6204; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_7757 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec_7_1_addr : _GEN_6205; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire  _GEN_7767 = next_reg_LevelVec_10_0_valid | _GEN_6207; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_7768 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec_7_0_addr : _GEN_6208; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] _GEN_7826 = next_reg_success_10 ? next_reg_finaladdr_7 : _GEN_5980; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 69:25]
  wire  _GEN_7828 = next_reg_success_10 ? _GEN_6216 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_7829 = next_reg_vmEnable_10 | _GEN_6201; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_7830 = next_reg_vmEnable_10 ? next_reg_LevelVec_7_2_addr : _GEN_6202; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_7832 = next_reg_vmEnable_10 ? _GEN_7756 : _GEN_6204; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_7833 = next_reg_vmEnable_10 ? _GEN_7757 : _GEN_6205; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_7835 = next_reg_vmEnable_10 ? _GEN_7767 : _GEN_6207; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_7836 = next_reg_vmEnable_10 ? _GEN_7768 : _GEN_6208; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_7842 = next_reg_vmEnable_10 ? _GEN_7826 : _next_reg_T_540; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22 74:23]
  wire  _GEN_7844 = next_reg_vmEnable_10 ? _GEN_7828 : _GEN_6216; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_7846 = 5'h1 == rd ? _next_reg_T_593 : _GEN_7695; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7847 = 5'h2 == rd ? _next_reg_T_593 : _GEN_7696; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7848 = 5'h3 == rd ? _next_reg_T_593 : _GEN_7697; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7849 = 5'h4 == rd ? _next_reg_T_593 : _GEN_7698; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7850 = 5'h5 == rd ? _next_reg_T_593 : _GEN_7699; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7851 = 5'h6 == rd ? _next_reg_T_593 : _GEN_7700; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7852 = 5'h7 == rd ? _next_reg_T_593 : _GEN_7701; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7853 = 5'h8 == rd ? _next_reg_T_593 : _GEN_7702; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7854 = 5'h9 == rd ? _next_reg_T_593 : _GEN_7703; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7855 = 5'ha == rd ? _next_reg_T_593 : _GEN_7704; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7856 = 5'hb == rd ? _next_reg_T_593 : _GEN_7705; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7857 = 5'hc == rd ? _next_reg_T_593 : _GEN_7706; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7858 = 5'hd == rd ? _next_reg_T_593 : _GEN_7707; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7859 = 5'he == rd ? _next_reg_T_593 : _GEN_7708; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7860 = 5'hf == rd ? _next_reg_T_593 : _GEN_7709; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7861 = 5'h10 == rd ? _next_reg_T_593 : _GEN_7710; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7862 = 5'h11 == rd ? _next_reg_T_593 : _GEN_7711; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7863 = 5'h12 == rd ? _next_reg_T_593 : _GEN_7712; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7864 = 5'h13 == rd ? _next_reg_T_593 : _GEN_7713; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7865 = 5'h14 == rd ? _next_reg_T_593 : _GEN_7714; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7866 = 5'h15 == rd ? _next_reg_T_593 : _GEN_7715; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7867 = 5'h16 == rd ? _next_reg_T_593 : _GEN_7716; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7868 = 5'h17 == rd ? _next_reg_T_593 : _GEN_7717; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7869 = 5'h18 == rd ? _next_reg_T_593 : _GEN_7718; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7870 = 5'h19 == rd ? _next_reg_T_593 : _GEN_7719; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7871 = 5'h1a == rd ? _next_reg_T_593 : _GEN_7720; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7872 = 5'h1b == rd ? _next_reg_T_593 : _GEN_7721; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7873 = 5'h1c == rd ? _next_reg_T_593 : _GEN_7722; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7874 = 5'h1d == rd ? _next_reg_T_593 : _GEN_7723; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7875 = 5'h1e == rd ? _next_reg_T_593 : _GEN_7724; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire [63:0] _GEN_7876 = 5'h1f == rd ? _next_reg_T_593 : _GEN_7725; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 270:{20,20}]
  wire  _GEN_7885 = _T_1308 | _GEN_5966; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 63:22]
  wire  _GEN_7886 = _T_1308 ? _GEN_7829 : _GEN_6201; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7887 = _T_1308 ? _GEN_7830 : _GEN_6202; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire  _GEN_7889 = _T_1308 ? _GEN_7832 : _GEN_6204; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7890 = _T_1308 ? _GEN_7833 : _GEN_6205; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire  _GEN_7892 = _T_1308 ? _GEN_7835 : _GEN_6207; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7893 = _T_1308 ? _GEN_7836 : _GEN_6208; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7899 = _T_1308 ? _GEN_7842 : _GEN_5980; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire  _GEN_7901 = _T_1308 ? _GEN_7844 : _GEN_6216; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [6:0] _GEN_7902 = _T_1308 ? 7'h40 : _GEN_5983; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 76:25]
  wire [63:0] _GEN_7904 = _T_1308 ? _GEN_7846 : _GEN_7695; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7905 = _T_1308 ? _GEN_7847 : _GEN_7696; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7906 = _T_1308 ? _GEN_7848 : _GEN_7697; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7907 = _T_1308 ? _GEN_7849 : _GEN_7698; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7908 = _T_1308 ? _GEN_7850 : _GEN_7699; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7909 = _T_1308 ? _GEN_7851 : _GEN_7700; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7910 = _T_1308 ? _GEN_7852 : _GEN_7701; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7911 = _T_1308 ? _GEN_7853 : _GEN_7702; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7912 = _T_1308 ? _GEN_7854 : _GEN_7703; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7913 = _T_1308 ? _GEN_7855 : _GEN_7704; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7914 = _T_1308 ? _GEN_7856 : _GEN_7705; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7915 = _T_1308 ? _GEN_7857 : _GEN_7706; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7916 = _T_1308 ? _GEN_7858 : _GEN_7707; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7917 = _T_1308 ? _GEN_7859 : _GEN_7708; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7918 = _T_1308 ? _GEN_7860 : _GEN_7709; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7919 = _T_1308 ? _GEN_7861 : _GEN_7710; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7920 = _T_1308 ? _GEN_7862 : _GEN_7711; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7921 = _T_1308 ? _GEN_7863 : _GEN_7712; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7922 = _T_1308 ? _GEN_7864 : _GEN_7713; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7923 = _T_1308 ? _GEN_7865 : _GEN_7714; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7924 = _T_1308 ? _GEN_7866 : _GEN_7715; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7925 = _T_1308 ? _GEN_7867 : _GEN_7716; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7926 = _T_1308 ? _GEN_7868 : _GEN_7717; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7927 = _T_1308 ? _GEN_7869 : _GEN_7718; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7928 = _T_1308 ? _GEN_7870 : _GEN_7719; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7929 = _T_1308 ? _GEN_7871 : _GEN_7720; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7930 = _T_1308 ? _GEN_7872 : _GEN_7721; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7931 = _T_1308 ? _GEN_7873 : _GEN_7722; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7932 = _T_1308 ? _GEN_7874 : _GEN_7723; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7933 = _T_1308 ? _GEN_7875 : _GEN_7724; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire [63:0] _GEN_7934 = _T_1308 ? _GEN_7876 : _GEN_7725; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 267:24]
  wire  _GEN_7958 = next_reg_LevelVec_10_1_valid | _GEN_7889; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_7959 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec_7_1_addr : _GEN_7890; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire  _GEN_7969 = next_reg_LevelVec_10_0_valid | _GEN_7892; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_7970 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec_7_0_addr : _GEN_7893; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] _GEN_8028 = success_8 ? finaladdr_5 : _GEN_6214; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 97:26]
  wire  _GEN_8030 = success_8 ? _GEN_7901 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_8031 = next_reg_vmEnable_10 | _GEN_7886; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_8032 = next_reg_vmEnable_10 ? next_reg_LevelVec_7_2_addr : _GEN_7887; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_8034 = next_reg_vmEnable_10 ? _GEN_7958 : _GEN_7889; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_8035 = next_reg_vmEnable_10 ? _GEN_7959 : _GEN_7890; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_8037 = next_reg_vmEnable_10 ? _GEN_7969 : _GEN_7892; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_8038 = next_reg_vmEnable_10 ? _GEN_7970 : _GEN_7893; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_8044 = next_reg_vmEnable_10 ? _GEN_8028 : _next_reg_T_540; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22 102:24]
  wire  _GEN_8046 = next_reg_vmEnable_10 ? _GEN_8030 : _GEN_7901; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_8053 = _T_1315 | _GEN_6200; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 92:23]
  wire  _GEN_8054 = _T_1315 ? _GEN_8031 : _GEN_7886; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24]
  wire [63:0] _GEN_8055 = _T_1315 ? _GEN_8032 : _GEN_7887; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24]
  wire  _GEN_8057 = _T_1315 ? _GEN_8034 : _GEN_7889; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24]
  wire [63:0] _GEN_8058 = _T_1315 ? _GEN_8035 : _GEN_7890; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24]
  wire  _GEN_8060 = _T_1315 ? _GEN_8037 : _GEN_7892; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24]
  wire [63:0] _GEN_8061 = _T_1315 ? _GEN_8038 : _GEN_7893; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24]
  wire [63:0] _GEN_8067 = _T_1315 ? _GEN_8044 : _GEN_6214; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24]
  wire  _GEN_8069 = _T_1315 ? _GEN_8046 : _GEN_7901; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24]
  wire [6:0] _GEN_8070 = _T_1315 ? 7'h40 : _GEN_6217; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 104:26]
  wire [63:0] _GEN_8071 = _T_1315 ? _GEN_910 : _GEN_6218; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 272:24 src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:26]
  wire  _GEN_8127 = next_reg_LevelVec_10_1_valid | _GEN_8057; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_8128 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec_8_1_addr : _GEN_8058; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire  _GEN_8138 = next_reg_LevelVec_10_0_valid | _GEN_8060; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_8139 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec_8_0_addr : _GEN_8061; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] _GEN_8197 = next_reg_success_10 ? next_reg_finaladdr_8 : _GEN_7899; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 69:25]
  wire  _GEN_8199 = next_reg_success_10 ? _GEN_8069 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 68:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_8200 = next_reg_vmEnable_10 | _GEN_8054; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_8201 = next_reg_vmEnable_10 ? next_reg_LevelVec_8_2_addr : _GEN_8055; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_8203 = next_reg_vmEnable_10 ? _GEN_8127 : _GEN_8057; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_8204 = next_reg_vmEnable_10 ? _GEN_8128 : _GEN_8058; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire  _GEN_8206 = next_reg_vmEnable_10 ? _GEN_8138 : _GEN_8060; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_8207 = next_reg_vmEnable_10 ? _GEN_8139 : _GEN_8061; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_8213 = next_reg_vmEnable_10 ? _GEN_8197 : _next_reg_T_601; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22 74:23]
  wire  _GEN_8215 = next_reg_vmEnable_10 ? _GEN_8199 : _GEN_8069; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 64:22]
  wire [63:0] _GEN_8217 = 5'h1 == _T_1012 ? _next_reg_T_654 : _GEN_7904; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8218 = 5'h2 == _T_1012 ? _next_reg_T_654 : _GEN_7905; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8219 = 5'h3 == _T_1012 ? _next_reg_T_654 : _GEN_7906; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8220 = 5'h4 == _T_1012 ? _next_reg_T_654 : _GEN_7907; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8221 = 5'h5 == _T_1012 ? _next_reg_T_654 : _GEN_7908; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8222 = 5'h6 == _T_1012 ? _next_reg_T_654 : _GEN_7909; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8223 = 5'h7 == _T_1012 ? _next_reg_T_654 : _GEN_7910; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8224 = 5'h8 == _T_1012 ? _next_reg_T_654 : _GEN_7911; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8225 = 5'h9 == _T_1012 ? _next_reg_T_654 : _GEN_7912; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8226 = 5'ha == _T_1012 ? _next_reg_T_654 : _GEN_7913; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8227 = 5'hb == _T_1012 ? _next_reg_T_654 : _GEN_7914; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8228 = 5'hc == _T_1012 ? _next_reg_T_654 : _GEN_7915; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8229 = 5'hd == _T_1012 ? _next_reg_T_654 : _GEN_7916; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8230 = 5'he == _T_1012 ? _next_reg_T_654 : _GEN_7917; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8231 = 5'hf == _T_1012 ? _next_reg_T_654 : _GEN_7918; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8232 = 5'h10 == _T_1012 ? _next_reg_T_654 : _GEN_7919; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8233 = 5'h11 == _T_1012 ? _next_reg_T_654 : _GEN_7920; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8234 = 5'h12 == _T_1012 ? _next_reg_T_654 : _GEN_7921; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8235 = 5'h13 == _T_1012 ? _next_reg_T_654 : _GEN_7922; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8236 = 5'h14 == _T_1012 ? _next_reg_T_654 : _GEN_7923; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8237 = 5'h15 == _T_1012 ? _next_reg_T_654 : _GEN_7924; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8238 = 5'h16 == _T_1012 ? _next_reg_T_654 : _GEN_7925; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8239 = 5'h17 == _T_1012 ? _next_reg_T_654 : _GEN_7926; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8240 = 5'h18 == _T_1012 ? _next_reg_T_654 : _GEN_7927; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8241 = 5'h19 == _T_1012 ? _next_reg_T_654 : _GEN_7928; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8242 = 5'h1a == _T_1012 ? _next_reg_T_654 : _GEN_7929; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8243 = 5'h1b == _T_1012 ? _next_reg_T_654 : _GEN_7930; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8244 = 5'h1c == _T_1012 ? _next_reg_T_654 : _GEN_7931; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8245 = 5'h1d == _T_1012 ? _next_reg_T_654 : _GEN_7932; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8246 = 5'h1e == _T_1012 ? _next_reg_T_654 : _GEN_7933; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire [63:0] _GEN_8247 = 5'h1f == _T_1012 ? _next_reg_T_654 : _GEN_7934; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 281:{28,28}]
  wire  _GEN_8256 = _T_1376 | _GEN_7885; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 63:22]
  wire  _GEN_8257 = _T_1376 ? _GEN_8200 : _GEN_8054; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8258 = _T_1376 ? _GEN_8201 : _GEN_8055; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire  _GEN_8260 = _T_1376 ? _GEN_8203 : _GEN_8057; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8261 = _T_1376 ? _GEN_8204 : _GEN_8058; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire  _GEN_8263 = _T_1376 ? _GEN_8206 : _GEN_8060; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8264 = _T_1376 ? _GEN_8207 : _GEN_8061; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8270 = _T_1376 ? _GEN_8213 : _GEN_7899; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire  _GEN_8272 = _T_1376 ? _GEN_8215 : _GEN_8069; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [6:0] _GEN_8273 = _T_1376 ? 7'h40 : _GEN_7902; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 76:25]
  wire [63:0] _GEN_8275 = _T_1376 ? _GEN_8217 : _GEN_7904; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8276 = _T_1376 ? _GEN_8218 : _GEN_7905; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8277 = _T_1376 ? _GEN_8219 : _GEN_7906; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8278 = _T_1376 ? _GEN_8220 : _GEN_7907; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8279 = _T_1376 ? _GEN_8221 : _GEN_7908; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8280 = _T_1376 ? _GEN_8222 : _GEN_7909; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8281 = _T_1376 ? _GEN_8223 : _GEN_7910; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8282 = _T_1376 ? _GEN_8224 : _GEN_7911; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8283 = _T_1376 ? _GEN_8225 : _GEN_7912; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8284 = _T_1376 ? _GEN_8226 : _GEN_7913; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8285 = _T_1376 ? _GEN_8227 : _GEN_7914; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8286 = _T_1376 ? _GEN_8228 : _GEN_7915; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8287 = _T_1376 ? _GEN_8229 : _GEN_7916; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8288 = _T_1376 ? _GEN_8230 : _GEN_7917; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8289 = _T_1376 ? _GEN_8231 : _GEN_7918; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8290 = _T_1376 ? _GEN_8232 : _GEN_7919; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8291 = _T_1376 ? _GEN_8233 : _GEN_7920; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8292 = _T_1376 ? _GEN_8234 : _GEN_7921; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8293 = _T_1376 ? _GEN_8235 : _GEN_7922; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8294 = _T_1376 ? _GEN_8236 : _GEN_7923; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8295 = _T_1376 ? _GEN_8237 : _GEN_7924; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8296 = _T_1376 ? _GEN_8238 : _GEN_7925; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8297 = _T_1376 ? _GEN_8239 : _GEN_7926; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8298 = _T_1376 ? _GEN_8240 : _GEN_7927; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8299 = _T_1376 ? _GEN_8241 : _GEN_7928; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8300 = _T_1376 ? _GEN_8242 : _GEN_7929; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8301 = _T_1376 ? _GEN_8243 : _GEN_7930; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8302 = _T_1376 ? _GEN_8244 : _GEN_7931; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8303 = _T_1376 ? _GEN_8245 : _GEN_7932; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8304 = _T_1376 ? _GEN_8246 : _GEN_7933; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire [63:0] _GEN_8305 = _T_1376 ? _GEN_8247 : _GEN_7934; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 278:22]
  wire  _GEN_8361 = next_reg_LevelVec_10_1_valid | _GEN_8260; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_8362 = next_reg_LevelVec_10_1_valid ? next_reg_LevelVec_8_1_addr : _GEN_8261; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire  _GEN_8372 = next_reg_LevelVec_10_0_valid | _GEN_8263; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 144:38 271:41]
  wire [63:0] _GEN_8373 = next_reg_LevelVec_10_0_valid ? next_reg_LevelVec_8_0_addr : _GEN_8264; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 145:38 271:41]
  wire [63:0] _GEN_8431 = success_8 ? finaladdr_6 : _GEN_8067; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 97:26]
  wire  _GEN_8433 = success_8 ? _GEN_8272 : 1'h1; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 96:23 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_8434 = next_reg_vmEnable_10 | _GEN_8257; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_8435 = next_reg_vmEnable_10 ? next_reg_LevelVec_8_2_addr : _GEN_8258; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_8437 = next_reg_vmEnable_10 ? _GEN_8361 : _GEN_8260; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_8438 = next_reg_vmEnable_10 ? _GEN_8362 : _GEN_8261; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_8440 = next_reg_vmEnable_10 ? _GEN_8372 : _GEN_8263; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_8441 = next_reg_vmEnable_10 ? _GEN_8373 : _GEN_8264; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire [63:0] _GEN_8447 = next_reg_vmEnable_10 ? _GEN_8431 : _next_reg_T_601; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22 102:24]
  wire  _GEN_8449 = next_reg_vmEnable_10 ? _GEN_8433 : _GEN_8272; // @[src/main/scala/rvspeccore/core/tool/LoadStore.scala 93:22]
  wire  _GEN_8490 = _T_1385 | _GEN_8053; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 92:23]
  wire  _GEN_8491 = _T_1385 ? _GEN_8434 : _GEN_8257; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22]
  wire [63:0] _GEN_8492 = _T_1385 ? _GEN_8435 : _GEN_8258; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22]
  wire  _GEN_8494 = _T_1385 ? _GEN_8437 : _GEN_8260; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22]
  wire [63:0] _GEN_8495 = _T_1385 ? _GEN_8438 : _GEN_8261; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22]
  wire  _GEN_8497 = _T_1385 ? _GEN_8440 : _GEN_8263; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22]
  wire [63:0] _GEN_8498 = _T_1385 ? _GEN_8441 : _GEN_8264; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22]
  wire [63:0] _GEN_8504 = _T_1385 ? _GEN_8447 : _GEN_8067; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22]
  wire  _GEN_8506 = _T_1385 ? _GEN_8449 : _GEN_8272; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22]
  wire [6:0] _GEN_8507 = _T_1385 ? 7'h40 : _GEN_8070; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 104:26]
  wire [63:0] _GEN_8508 = _T_1385 ? _GEN_6191 : _GEN_8071; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 283:22 src/main/scala/rvspeccore/core/tool/LoadStore.scala 105:26]
  wire [63:0] _next_reg_T_811 = _GEN_6513 + imm; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:44]
  wire  next_reg_signBit_17 = _next_reg_T_811[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_814 = next_reg_signBit_17 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_815 = {_next_reg_T_814,_next_reg_T_811[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_8510 = 5'h1 == rd ? _next_reg_T_815 : _GEN_8275; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8511 = 5'h2 == rd ? _next_reg_T_815 : _GEN_8276; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8512 = 5'h3 == rd ? _next_reg_T_815 : _GEN_8277; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8513 = 5'h4 == rd ? _next_reg_T_815 : _GEN_8278; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8514 = 5'h5 == rd ? _next_reg_T_815 : _GEN_8279; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8515 = 5'h6 == rd ? _next_reg_T_815 : _GEN_8280; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8516 = 5'h7 == rd ? _next_reg_T_815 : _GEN_8281; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8517 = 5'h8 == rd ? _next_reg_T_815 : _GEN_8282; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8518 = 5'h9 == rd ? _next_reg_T_815 : _GEN_8283; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8519 = 5'ha == rd ? _next_reg_T_815 : _GEN_8284; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8520 = 5'hb == rd ? _next_reg_T_815 : _GEN_8285; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8521 = 5'hc == rd ? _next_reg_T_815 : _GEN_8286; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8522 = 5'hd == rd ? _next_reg_T_815 : _GEN_8287; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8523 = 5'he == rd ? _next_reg_T_815 : _GEN_8288; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8524 = 5'hf == rd ? _next_reg_T_815 : _GEN_8289; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8525 = 5'h10 == rd ? _next_reg_T_815 : _GEN_8290; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8526 = 5'h11 == rd ? _next_reg_T_815 : _GEN_8291; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8527 = 5'h12 == rd ? _next_reg_T_815 : _GEN_8292; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8528 = 5'h13 == rd ? _next_reg_T_815 : _GEN_8293; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8529 = 5'h14 == rd ? _next_reg_T_815 : _GEN_8294; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8530 = 5'h15 == rd ? _next_reg_T_815 : _GEN_8295; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8531 = 5'h16 == rd ? _next_reg_T_815 : _GEN_8296; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8532 = 5'h17 == rd ? _next_reg_T_815 : _GEN_8297; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8533 = 5'h18 == rd ? _next_reg_T_815 : _GEN_8298; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8534 = 5'h19 == rd ? _next_reg_T_815 : _GEN_8299; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8535 = 5'h1a == rd ? _next_reg_T_815 : _GEN_8300; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8536 = 5'h1b == rd ? _next_reg_T_815 : _GEN_8301; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8537 = 5'h1c == rd ? _next_reg_T_815 : _GEN_8302; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8538 = 5'h1d == rd ? _next_reg_T_815 : _GEN_8303; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8539 = 5'h1e == rd ? _next_reg_T_815 : _GEN_8304; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8540 = 5'h1f == rd ? _next_reg_T_815 : _GEN_8305; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 293:{20,20}]
  wire [63:0] _GEN_8550 = _T_1452 ? _GEN_8510 : _GEN_8275; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8551 = _T_1452 ? _GEN_8511 : _GEN_8276; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8552 = _T_1452 ? _GEN_8512 : _GEN_8277; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8553 = _T_1452 ? _GEN_8513 : _GEN_8278; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8554 = _T_1452 ? _GEN_8514 : _GEN_8279; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8555 = _T_1452 ? _GEN_8515 : _GEN_8280; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8556 = _T_1452 ? _GEN_8516 : _GEN_8281; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8557 = _T_1452 ? _GEN_8517 : _GEN_8282; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8558 = _T_1452 ? _GEN_8518 : _GEN_8283; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8559 = _T_1452 ? _GEN_8519 : _GEN_8284; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8560 = _T_1452 ? _GEN_8520 : _GEN_8285; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8561 = _T_1452 ? _GEN_8521 : _GEN_8286; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8562 = _T_1452 ? _GEN_8522 : _GEN_8287; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8563 = _T_1452 ? _GEN_8523 : _GEN_8288; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8564 = _T_1452 ? _GEN_8524 : _GEN_8289; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8565 = _T_1452 ? _GEN_8525 : _GEN_8290; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8566 = _T_1452 ? _GEN_8526 : _GEN_8291; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8567 = _T_1452 ? _GEN_8527 : _GEN_8292; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8568 = _T_1452 ? _GEN_8528 : _GEN_8293; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8569 = _T_1452 ? _GEN_8529 : _GEN_8294; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8570 = _T_1452 ? _GEN_8530 : _GEN_8295; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8571 = _T_1452 ? _GEN_8531 : _GEN_8296; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8572 = _T_1452 ? _GEN_8532 : _GEN_8297; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8573 = _T_1452 ? _GEN_8533 : _GEN_8298; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8574 = _T_1452 ? _GEN_8534 : _GEN_8299; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8575 = _T_1452 ? _GEN_8535 : _GEN_8300; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8576 = _T_1452 ? _GEN_8536 : _GEN_8301; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8577 = _T_1452 ? _GEN_8537 : _GEN_8302; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8578 = _T_1452 ? _GEN_8538 : _GEN_8303; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8579 = _T_1452 ? _GEN_8539 : _GEN_8304; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [63:0] _GEN_8580 = _T_1452 ? _GEN_8540 : _GEN_8305; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 290:25]
  wire [31:0] _next_reg_T_821 = _GEN_6765[31:0] + _GEN_6191[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:66]
  wire  next_reg_signBit_18 = _next_reg_T_821[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_823 = next_reg_signBit_18 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_824 = {_next_reg_T_823,_next_reg_T_821}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_8646 = 5'h1 == _T_1012 ? _next_reg_T_824 : _GEN_8550; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8647 = 5'h2 == _T_1012 ? _next_reg_T_824 : _GEN_8551; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8648 = 5'h3 == _T_1012 ? _next_reg_T_824 : _GEN_8552; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8649 = 5'h4 == _T_1012 ? _next_reg_T_824 : _GEN_8553; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8650 = 5'h5 == _T_1012 ? _next_reg_T_824 : _GEN_8554; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8651 = 5'h6 == _T_1012 ? _next_reg_T_824 : _GEN_8555; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8652 = 5'h7 == _T_1012 ? _next_reg_T_824 : _GEN_8556; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8653 = 5'h8 == _T_1012 ? _next_reg_T_824 : _GEN_8557; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8654 = 5'h9 == _T_1012 ? _next_reg_T_824 : _GEN_8558; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8655 = 5'ha == _T_1012 ? _next_reg_T_824 : _GEN_8559; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8656 = 5'hb == _T_1012 ? _next_reg_T_824 : _GEN_8560; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8657 = 5'hc == _T_1012 ? _next_reg_T_824 : _GEN_8561; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8658 = 5'hd == _T_1012 ? _next_reg_T_824 : _GEN_8562; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8659 = 5'he == _T_1012 ? _next_reg_T_824 : _GEN_8563; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8660 = 5'hf == _T_1012 ? _next_reg_T_824 : _GEN_8564; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8661 = 5'h10 == _T_1012 ? _next_reg_T_824 : _GEN_8565; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8662 = 5'h11 == _T_1012 ? _next_reg_T_824 : _GEN_8566; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8663 = 5'h12 == _T_1012 ? _next_reg_T_824 : _GEN_8567; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8664 = 5'h13 == _T_1012 ? _next_reg_T_824 : _GEN_8568; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8665 = 5'h14 == _T_1012 ? _next_reg_T_824 : _GEN_8569; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8666 = 5'h15 == _T_1012 ? _next_reg_T_824 : _GEN_8570; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8667 = 5'h16 == _T_1012 ? _next_reg_T_824 : _GEN_8571; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8668 = 5'h17 == _T_1012 ? _next_reg_T_824 : _GEN_8572; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8669 = 5'h18 == _T_1012 ? _next_reg_T_824 : _GEN_8573; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8670 = 5'h19 == _T_1012 ? _next_reg_T_824 : _GEN_8574; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8671 = 5'h1a == _T_1012 ? _next_reg_T_824 : _GEN_8575; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8672 = 5'h1b == _T_1012 ? _next_reg_T_824 : _GEN_8576; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8673 = 5'h1c == _T_1012 ? _next_reg_T_824 : _GEN_8577; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8674 = 5'h1d == _T_1012 ? _next_reg_T_824 : _GEN_8578; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8675 = 5'h1e == _T_1012 ? _next_reg_T_824 : _GEN_8579; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8676 = 5'h1f == _T_1012 ? _next_reg_T_824 : _GEN_8580; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 299:{28,28}]
  wire [63:0] _GEN_8685 = _T_1459 ? _GEN_8646 : _GEN_8550; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8686 = _T_1459 ? _GEN_8647 : _GEN_8551; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8687 = _T_1459 ? _GEN_8648 : _GEN_8552; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8688 = _T_1459 ? _GEN_8649 : _GEN_8553; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8689 = _T_1459 ? _GEN_8650 : _GEN_8554; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8690 = _T_1459 ? _GEN_8651 : _GEN_8555; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8691 = _T_1459 ? _GEN_8652 : _GEN_8556; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8692 = _T_1459 ? _GEN_8653 : _GEN_8557; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8693 = _T_1459 ? _GEN_8654 : _GEN_8558; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8694 = _T_1459 ? _GEN_8655 : _GEN_8559; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8695 = _T_1459 ? _GEN_8656 : _GEN_8560; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8696 = _T_1459 ? _GEN_8657 : _GEN_8561; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8697 = _T_1459 ? _GEN_8658 : _GEN_8562; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8698 = _T_1459 ? _GEN_8659 : _GEN_8563; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8699 = _T_1459 ? _GEN_8660 : _GEN_8564; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8700 = _T_1459 ? _GEN_8661 : _GEN_8565; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8701 = _T_1459 ? _GEN_8662 : _GEN_8566; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8702 = _T_1459 ? _GEN_8663 : _GEN_8567; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8703 = _T_1459 ? _GEN_8664 : _GEN_8568; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8704 = _T_1459 ? _GEN_8665 : _GEN_8569; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8705 = _T_1459 ? _GEN_8666 : _GEN_8570; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8706 = _T_1459 ? _GEN_8667 : _GEN_8571; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8707 = _T_1459 ? _GEN_8668 : _GEN_8572; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8708 = _T_1459 ? _GEN_8669 : _GEN_8573; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8709 = _T_1459 ? _GEN_8670 : _GEN_8574; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8710 = _T_1459 ? _GEN_8671 : _GEN_8575; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8711 = _T_1459 ? _GEN_8672 : _GEN_8576; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8712 = _T_1459 ? _GEN_8673 : _GEN_8577; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8713 = _T_1459 ? _GEN_8674 : _GEN_8578; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8714 = _T_1459 ? _GEN_8675 : _GEN_8579; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [63:0] _GEN_8715 = _T_1459 ? _GEN_8676 : _GEN_8580; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 297:24]
  wire [31:0] _next_reg_T_830 = _GEN_6765[31:0] - _GEN_6191[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:66]
  wire  next_reg_signBit_19 = _next_reg_T_830[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_832 = next_reg_signBit_19 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_833 = {_next_reg_T_832,_next_reg_T_830}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_8781 = 5'h1 == _T_1012 ? _next_reg_T_833 : _GEN_8685; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8782 = 5'h2 == _T_1012 ? _next_reg_T_833 : _GEN_8686; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8783 = 5'h3 == _T_1012 ? _next_reg_T_833 : _GEN_8687; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8784 = 5'h4 == _T_1012 ? _next_reg_T_833 : _GEN_8688; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8785 = 5'h5 == _T_1012 ? _next_reg_T_833 : _GEN_8689; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8786 = 5'h6 == _T_1012 ? _next_reg_T_833 : _GEN_8690; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8787 = 5'h7 == _T_1012 ? _next_reg_T_833 : _GEN_8691; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8788 = 5'h8 == _T_1012 ? _next_reg_T_833 : _GEN_8692; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8789 = 5'h9 == _T_1012 ? _next_reg_T_833 : _GEN_8693; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8790 = 5'ha == _T_1012 ? _next_reg_T_833 : _GEN_8694; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8791 = 5'hb == _T_1012 ? _next_reg_T_833 : _GEN_8695; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8792 = 5'hc == _T_1012 ? _next_reg_T_833 : _GEN_8696; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8793 = 5'hd == _T_1012 ? _next_reg_T_833 : _GEN_8697; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8794 = 5'he == _T_1012 ? _next_reg_T_833 : _GEN_8698; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8795 = 5'hf == _T_1012 ? _next_reg_T_833 : _GEN_8699; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8796 = 5'h10 == _T_1012 ? _next_reg_T_833 : _GEN_8700; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8797 = 5'h11 == _T_1012 ? _next_reg_T_833 : _GEN_8701; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8798 = 5'h12 == _T_1012 ? _next_reg_T_833 : _GEN_8702; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8799 = 5'h13 == _T_1012 ? _next_reg_T_833 : _GEN_8703; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8800 = 5'h14 == _T_1012 ? _next_reg_T_833 : _GEN_8704; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8801 = 5'h15 == _T_1012 ? _next_reg_T_833 : _GEN_8705; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8802 = 5'h16 == _T_1012 ? _next_reg_T_833 : _GEN_8706; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8803 = 5'h17 == _T_1012 ? _next_reg_T_833 : _GEN_8707; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8804 = 5'h18 == _T_1012 ? _next_reg_T_833 : _GEN_8708; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8805 = 5'h19 == _T_1012 ? _next_reg_T_833 : _GEN_8709; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8806 = 5'h1a == _T_1012 ? _next_reg_T_833 : _GEN_8710; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8807 = 5'h1b == _T_1012 ? _next_reg_T_833 : _GEN_8711; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8808 = 5'h1c == _T_1012 ? _next_reg_T_833 : _GEN_8712; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8809 = 5'h1d == _T_1012 ? _next_reg_T_833 : _GEN_8713; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8810 = 5'h1e == _T_1012 ? _next_reg_T_833 : _GEN_8714; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8811 = 5'h1f == _T_1012 ? _next_reg_T_833 : _GEN_8715; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 303:{28,28}]
  wire [63:0] _GEN_8820 = _T_1467 ? _GEN_8781 : _GEN_8685; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8821 = _T_1467 ? _GEN_8782 : _GEN_8686; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8822 = _T_1467 ? _GEN_8783 : _GEN_8687; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8823 = _T_1467 ? _GEN_8784 : _GEN_8688; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8824 = _T_1467 ? _GEN_8785 : _GEN_8689; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8825 = _T_1467 ? _GEN_8786 : _GEN_8690; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8826 = _T_1467 ? _GEN_8787 : _GEN_8691; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8827 = _T_1467 ? _GEN_8788 : _GEN_8692; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8828 = _T_1467 ? _GEN_8789 : _GEN_8693; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8829 = _T_1467 ? _GEN_8790 : _GEN_8694; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8830 = _T_1467 ? _GEN_8791 : _GEN_8695; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8831 = _T_1467 ? _GEN_8792 : _GEN_8696; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8832 = _T_1467 ? _GEN_8793 : _GEN_8697; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8833 = _T_1467 ? _GEN_8794 : _GEN_8698; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8834 = _T_1467 ? _GEN_8795 : _GEN_8699; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8835 = _T_1467 ? _GEN_8796 : _GEN_8700; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8836 = _T_1467 ? _GEN_8797 : _GEN_8701; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8837 = _T_1467 ? _GEN_8798 : _GEN_8702; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8838 = _T_1467 ? _GEN_8799 : _GEN_8703; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8839 = _T_1467 ? _GEN_8800 : _GEN_8704; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8840 = _T_1467 ? _GEN_8801 : _GEN_8705; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8841 = _T_1467 ? _GEN_8802 : _GEN_8706; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8842 = _T_1467 ? _GEN_8803 : _GEN_8707; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8843 = _T_1467 ? _GEN_8804 : _GEN_8708; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8844 = _T_1467 ? _GEN_8805 : _GEN_8709; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8845 = _T_1467 ? _GEN_8806 : _GEN_8710; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8846 = _T_1467 ? _GEN_8807 : _GEN_8711; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8847 = _T_1467 ? _GEN_8808 : _GEN_8712; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8848 = _T_1467 ? _GEN_8809 : _GEN_8713; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8849 = _T_1467 ? _GEN_8810 : _GEN_8714; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [63:0] _GEN_8850 = _T_1467 ? _GEN_8811 : _GEN_8715; // @[src/main/scala/rvspeccore/core/spec/instset/CExtension.scala 301:24]
  wire [127:0] _next_reg_T_834 = _GEN_101 * _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:65]
  wire [63:0] _GEN_8852 = 5'h1 == rd ? _next_reg_T_834[63:0] : _GEN_8820; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8853 = 5'h2 == rd ? _next_reg_T_834[63:0] : _GEN_8821; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8854 = 5'h3 == rd ? _next_reg_T_834[63:0] : _GEN_8822; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8855 = 5'h4 == rd ? _next_reg_T_834[63:0] : _GEN_8823; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8856 = 5'h5 == rd ? _next_reg_T_834[63:0] : _GEN_8824; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8857 = 5'h6 == rd ? _next_reg_T_834[63:0] : _GEN_8825; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8858 = 5'h7 == rd ? _next_reg_T_834[63:0] : _GEN_8826; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8859 = 5'h8 == rd ? _next_reg_T_834[63:0] : _GEN_8827; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8860 = 5'h9 == rd ? _next_reg_T_834[63:0] : _GEN_8828; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8861 = 5'ha == rd ? _next_reg_T_834[63:0] : _GEN_8829; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8862 = 5'hb == rd ? _next_reg_T_834[63:0] : _GEN_8830; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8863 = 5'hc == rd ? _next_reg_T_834[63:0] : _GEN_8831; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8864 = 5'hd == rd ? _next_reg_T_834[63:0] : _GEN_8832; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8865 = 5'he == rd ? _next_reg_T_834[63:0] : _GEN_8833; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8866 = 5'hf == rd ? _next_reg_T_834[63:0] : _GEN_8834; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8867 = 5'h10 == rd ? _next_reg_T_834[63:0] : _GEN_8835; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8868 = 5'h11 == rd ? _next_reg_T_834[63:0] : _GEN_8836; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8869 = 5'h12 == rd ? _next_reg_T_834[63:0] : _GEN_8837; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8870 = 5'h13 == rd ? _next_reg_T_834[63:0] : _GEN_8838; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8871 = 5'h14 == rd ? _next_reg_T_834[63:0] : _GEN_8839; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8872 = 5'h15 == rd ? _next_reg_T_834[63:0] : _GEN_8840; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8873 = 5'h16 == rd ? _next_reg_T_834[63:0] : _GEN_8841; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8874 = 5'h17 == rd ? _next_reg_T_834[63:0] : _GEN_8842; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8875 = 5'h18 == rd ? _next_reg_T_834[63:0] : _GEN_8843; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8876 = 5'h19 == rd ? _next_reg_T_834[63:0] : _GEN_8844; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8877 = 5'h1a == rd ? _next_reg_T_834[63:0] : _GEN_8845; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8878 = 5'h1b == rd ? _next_reg_T_834[63:0] : _GEN_8846; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8879 = 5'h1c == rd ? _next_reg_T_834[63:0] : _GEN_8847; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8880 = 5'h1d == rd ? _next_reg_T_834[63:0] : _GEN_8848; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8881 = 5'h1e == rd ? _next_reg_T_834[63:0] : _GEN_8849; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8882 = 5'h1f == rd ? _next_reg_T_834[63:0] : _GEN_8850; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:{48,48}]
  wire [63:0] _GEN_8891 = _T_1475 ? _GEN_8852 : _GEN_8820; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8892 = _T_1475 ? _GEN_8853 : _GEN_8821; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8893 = _T_1475 ? _GEN_8854 : _GEN_8822; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8894 = _T_1475 ? _GEN_8855 : _GEN_8823; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8895 = _T_1475 ? _GEN_8856 : _GEN_8824; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8896 = _T_1475 ? _GEN_8857 : _GEN_8825; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8897 = _T_1475 ? _GEN_8858 : _GEN_8826; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8898 = _T_1475 ? _GEN_8859 : _GEN_8827; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8899 = _T_1475 ? _GEN_8860 : _GEN_8828; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8900 = _T_1475 ? _GEN_8861 : _GEN_8829; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8901 = _T_1475 ? _GEN_8862 : _GEN_8830; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8902 = _T_1475 ? _GEN_8863 : _GEN_8831; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8903 = _T_1475 ? _GEN_8864 : _GEN_8832; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8904 = _T_1475 ? _GEN_8865 : _GEN_8833; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8905 = _T_1475 ? _GEN_8866 : _GEN_8834; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8906 = _T_1475 ? _GEN_8867 : _GEN_8835; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8907 = _T_1475 ? _GEN_8868 : _GEN_8836; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8908 = _T_1475 ? _GEN_8869 : _GEN_8837; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8909 = _T_1475 ? _GEN_8870 : _GEN_8838; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8910 = _T_1475 ? _GEN_8871 : _GEN_8839; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8911 = _T_1475 ? _GEN_8872 : _GEN_8840; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8912 = _T_1475 ? _GEN_8873 : _GEN_8841; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8913 = _T_1475 ? _GEN_8874 : _GEN_8842; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8914 = _T_1475 ? _GEN_8875 : _GEN_8843; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8915 = _T_1475 ? _GEN_8876 : _GEN_8844; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8916 = _T_1475 ? _GEN_8877 : _GEN_8845; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8917 = _T_1475 ? _GEN_8878 : _GEN_8846; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8918 = _T_1475 ? _GEN_8879 : _GEN_8847; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8919 = _T_1475 ? _GEN_8880 : _GEN_8848; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8920 = _T_1475 ? _GEN_8881 : _GEN_8849; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [63:0] _GEN_8921 = _T_1475 ? _GEN_8882 : _GEN_8850; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 85:24]
  wire [127:0] _next_reg_T_839 = $signed(_T_325) * $signed(_T_326); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:95]
  wire [63:0] _GEN_8923 = 5'h1 == rd ? _next_reg_T_839[127:64] : _GEN_8891; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8924 = 5'h2 == rd ? _next_reg_T_839[127:64] : _GEN_8892; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8925 = 5'h3 == rd ? _next_reg_T_839[127:64] : _GEN_8893; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8926 = 5'h4 == rd ? _next_reg_T_839[127:64] : _GEN_8894; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8927 = 5'h5 == rd ? _next_reg_T_839[127:64] : _GEN_8895; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8928 = 5'h6 == rd ? _next_reg_T_839[127:64] : _GEN_8896; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8929 = 5'h7 == rd ? _next_reg_T_839[127:64] : _GEN_8897; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8930 = 5'h8 == rd ? _next_reg_T_839[127:64] : _GEN_8898; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8931 = 5'h9 == rd ? _next_reg_T_839[127:64] : _GEN_8899; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8932 = 5'ha == rd ? _next_reg_T_839[127:64] : _GEN_8900; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8933 = 5'hb == rd ? _next_reg_T_839[127:64] : _GEN_8901; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8934 = 5'hc == rd ? _next_reg_T_839[127:64] : _GEN_8902; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8935 = 5'hd == rd ? _next_reg_T_839[127:64] : _GEN_8903; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8936 = 5'he == rd ? _next_reg_T_839[127:64] : _GEN_8904; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8937 = 5'hf == rd ? _next_reg_T_839[127:64] : _GEN_8905; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8938 = 5'h10 == rd ? _next_reg_T_839[127:64] : _GEN_8906; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8939 = 5'h11 == rd ? _next_reg_T_839[127:64] : _GEN_8907; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8940 = 5'h12 == rd ? _next_reg_T_839[127:64] : _GEN_8908; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8941 = 5'h13 == rd ? _next_reg_T_839[127:64] : _GEN_8909; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8942 = 5'h14 == rd ? _next_reg_T_839[127:64] : _GEN_8910; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8943 = 5'h15 == rd ? _next_reg_T_839[127:64] : _GEN_8911; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8944 = 5'h16 == rd ? _next_reg_T_839[127:64] : _GEN_8912; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8945 = 5'h17 == rd ? _next_reg_T_839[127:64] : _GEN_8913; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8946 = 5'h18 == rd ? _next_reg_T_839[127:64] : _GEN_8914; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8947 = 5'h19 == rd ? _next_reg_T_839[127:64] : _GEN_8915; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8948 = 5'h1a == rd ? _next_reg_T_839[127:64] : _GEN_8916; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8949 = 5'h1b == rd ? _next_reg_T_839[127:64] : _GEN_8917; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8950 = 5'h1c == rd ? _next_reg_T_839[127:64] : _GEN_8918; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8951 = 5'h1d == rd ? _next_reg_T_839[127:64] : _GEN_8919; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8952 = 5'h1e == rd ? _next_reg_T_839[127:64] : _GEN_8920; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8953 = 5'h1f == rd ? _next_reg_T_839[127:64] : _GEN_8921; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:{48,48}]
  wire [63:0] _GEN_8962 = _T_1482 ? _GEN_8923 : _GEN_8891; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8963 = _T_1482 ? _GEN_8924 : _GEN_8892; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8964 = _T_1482 ? _GEN_8925 : _GEN_8893; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8965 = _T_1482 ? _GEN_8926 : _GEN_8894; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8966 = _T_1482 ? _GEN_8927 : _GEN_8895; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8967 = _T_1482 ? _GEN_8928 : _GEN_8896; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8968 = _T_1482 ? _GEN_8929 : _GEN_8897; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8969 = _T_1482 ? _GEN_8930 : _GEN_8898; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8970 = _T_1482 ? _GEN_8931 : _GEN_8899; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8971 = _T_1482 ? _GEN_8932 : _GEN_8900; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8972 = _T_1482 ? _GEN_8933 : _GEN_8901; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8973 = _T_1482 ? _GEN_8934 : _GEN_8902; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8974 = _T_1482 ? _GEN_8935 : _GEN_8903; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8975 = _T_1482 ? _GEN_8936 : _GEN_8904; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8976 = _T_1482 ? _GEN_8937 : _GEN_8905; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8977 = _T_1482 ? _GEN_8938 : _GEN_8906; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8978 = _T_1482 ? _GEN_8939 : _GEN_8907; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8979 = _T_1482 ? _GEN_8940 : _GEN_8908; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8980 = _T_1482 ? _GEN_8941 : _GEN_8909; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8981 = _T_1482 ? _GEN_8942 : _GEN_8910; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8982 = _T_1482 ? _GEN_8943 : _GEN_8911; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8983 = _T_1482 ? _GEN_8944 : _GEN_8912; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8984 = _T_1482 ? _GEN_8945 : _GEN_8913; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8985 = _T_1482 ? _GEN_8946 : _GEN_8914; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8986 = _T_1482 ? _GEN_8947 : _GEN_8915; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8987 = _T_1482 ? _GEN_8948 : _GEN_8916; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8988 = _T_1482 ? _GEN_8949 : _GEN_8917; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8989 = _T_1482 ? _GEN_8950 : _GEN_8918; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8990 = _T_1482 ? _GEN_8951 : _GEN_8919; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8991 = _T_1482 ? _GEN_8952 : _GEN_8920; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [63:0] _GEN_8992 = _T_1482 ? _GEN_8953 : _GEN_8921; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 86:24]
  wire [64:0] _next_reg_T_842 = {1'b0,$signed(_GEN_910)}; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:72]
  wire [128:0] _next_reg_T_843 = $signed(_T_325) * $signed(_next_reg_T_842); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:72]
  wire [127:0] _next_reg_T_846 = _next_reg_T_843[127:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:88]
  wire [63:0] _GEN_8994 = 5'h1 == rd ? _next_reg_T_846[127:64] : _GEN_8962; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_8995 = 5'h2 == rd ? _next_reg_T_846[127:64] : _GEN_8963; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_8996 = 5'h3 == rd ? _next_reg_T_846[127:64] : _GEN_8964; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_8997 = 5'h4 == rd ? _next_reg_T_846[127:64] : _GEN_8965; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_8998 = 5'h5 == rd ? _next_reg_T_846[127:64] : _GEN_8966; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_8999 = 5'h6 == rd ? _next_reg_T_846[127:64] : _GEN_8967; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9000 = 5'h7 == rd ? _next_reg_T_846[127:64] : _GEN_8968; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9001 = 5'h8 == rd ? _next_reg_T_846[127:64] : _GEN_8969; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9002 = 5'h9 == rd ? _next_reg_T_846[127:64] : _GEN_8970; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9003 = 5'ha == rd ? _next_reg_T_846[127:64] : _GEN_8971; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9004 = 5'hb == rd ? _next_reg_T_846[127:64] : _GEN_8972; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9005 = 5'hc == rd ? _next_reg_T_846[127:64] : _GEN_8973; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9006 = 5'hd == rd ? _next_reg_T_846[127:64] : _GEN_8974; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9007 = 5'he == rd ? _next_reg_T_846[127:64] : _GEN_8975; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9008 = 5'hf == rd ? _next_reg_T_846[127:64] : _GEN_8976; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9009 = 5'h10 == rd ? _next_reg_T_846[127:64] : _GEN_8977; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9010 = 5'h11 == rd ? _next_reg_T_846[127:64] : _GEN_8978; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9011 = 5'h12 == rd ? _next_reg_T_846[127:64] : _GEN_8979; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9012 = 5'h13 == rd ? _next_reg_T_846[127:64] : _GEN_8980; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9013 = 5'h14 == rd ? _next_reg_T_846[127:64] : _GEN_8981; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9014 = 5'h15 == rd ? _next_reg_T_846[127:64] : _GEN_8982; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9015 = 5'h16 == rd ? _next_reg_T_846[127:64] : _GEN_8983; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9016 = 5'h17 == rd ? _next_reg_T_846[127:64] : _GEN_8984; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9017 = 5'h18 == rd ? _next_reg_T_846[127:64] : _GEN_8985; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9018 = 5'h19 == rd ? _next_reg_T_846[127:64] : _GEN_8986; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9019 = 5'h1a == rd ? _next_reg_T_846[127:64] : _GEN_8987; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9020 = 5'h1b == rd ? _next_reg_T_846[127:64] : _GEN_8988; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9021 = 5'h1c == rd ? _next_reg_T_846[127:64] : _GEN_8989; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9022 = 5'h1d == rd ? _next_reg_T_846[127:64] : _GEN_8990; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9023 = 5'h1e == rd ? _next_reg_T_846[127:64] : _GEN_8991; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9024 = 5'h1f == rd ? _next_reg_T_846[127:64] : _GEN_8992; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:{48,48}]
  wire [63:0] _GEN_9033 = _T_1489 ? _GEN_8994 : _GEN_8962; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9034 = _T_1489 ? _GEN_8995 : _GEN_8963; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9035 = _T_1489 ? _GEN_8996 : _GEN_8964; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9036 = _T_1489 ? _GEN_8997 : _GEN_8965; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9037 = _T_1489 ? _GEN_8998 : _GEN_8966; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9038 = _T_1489 ? _GEN_8999 : _GEN_8967; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9039 = _T_1489 ? _GEN_9000 : _GEN_8968; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9040 = _T_1489 ? _GEN_9001 : _GEN_8969; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9041 = _T_1489 ? _GEN_9002 : _GEN_8970; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9042 = _T_1489 ? _GEN_9003 : _GEN_8971; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9043 = _T_1489 ? _GEN_9004 : _GEN_8972; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9044 = _T_1489 ? _GEN_9005 : _GEN_8973; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9045 = _T_1489 ? _GEN_9006 : _GEN_8974; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9046 = _T_1489 ? _GEN_9007 : _GEN_8975; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9047 = _T_1489 ? _GEN_9008 : _GEN_8976; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9048 = _T_1489 ? _GEN_9009 : _GEN_8977; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9049 = _T_1489 ? _GEN_9010 : _GEN_8978; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9050 = _T_1489 ? _GEN_9011 : _GEN_8979; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9051 = _T_1489 ? _GEN_9012 : _GEN_8980; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9052 = _T_1489 ? _GEN_9013 : _GEN_8981; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9053 = _T_1489 ? _GEN_9014 : _GEN_8982; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9054 = _T_1489 ? _GEN_9015 : _GEN_8983; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9055 = _T_1489 ? _GEN_9016 : _GEN_8984; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9056 = _T_1489 ? _GEN_9017 : _GEN_8985; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9057 = _T_1489 ? _GEN_9018 : _GEN_8986; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9058 = _T_1489 ? _GEN_9019 : _GEN_8987; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9059 = _T_1489 ? _GEN_9020 : _GEN_8988; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9060 = _T_1489 ? _GEN_9021 : _GEN_8989; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9061 = _T_1489 ? _GEN_9022 : _GEN_8990; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9062 = _T_1489 ? _GEN_9023 : _GEN_8991; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9063 = _T_1489 ? _GEN_9024 : _GEN_8992; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 87:24]
  wire [63:0] _GEN_9065 = 5'h1 == rd ? _next_reg_T_834[127:64] : _GEN_9033; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9066 = 5'h2 == rd ? _next_reg_T_834[127:64] : _GEN_9034; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9067 = 5'h3 == rd ? _next_reg_T_834[127:64] : _GEN_9035; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9068 = 5'h4 == rd ? _next_reg_T_834[127:64] : _GEN_9036; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9069 = 5'h5 == rd ? _next_reg_T_834[127:64] : _GEN_9037; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9070 = 5'h6 == rd ? _next_reg_T_834[127:64] : _GEN_9038; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9071 = 5'h7 == rd ? _next_reg_T_834[127:64] : _GEN_9039; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9072 = 5'h8 == rd ? _next_reg_T_834[127:64] : _GEN_9040; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9073 = 5'h9 == rd ? _next_reg_T_834[127:64] : _GEN_9041; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9074 = 5'ha == rd ? _next_reg_T_834[127:64] : _GEN_9042; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9075 = 5'hb == rd ? _next_reg_T_834[127:64] : _GEN_9043; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9076 = 5'hc == rd ? _next_reg_T_834[127:64] : _GEN_9044; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9077 = 5'hd == rd ? _next_reg_T_834[127:64] : _GEN_9045; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9078 = 5'he == rd ? _next_reg_T_834[127:64] : _GEN_9046; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9079 = 5'hf == rd ? _next_reg_T_834[127:64] : _GEN_9047; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9080 = 5'h10 == rd ? _next_reg_T_834[127:64] : _GEN_9048; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9081 = 5'h11 == rd ? _next_reg_T_834[127:64] : _GEN_9049; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9082 = 5'h12 == rd ? _next_reg_T_834[127:64] : _GEN_9050; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9083 = 5'h13 == rd ? _next_reg_T_834[127:64] : _GEN_9051; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9084 = 5'h14 == rd ? _next_reg_T_834[127:64] : _GEN_9052; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9085 = 5'h15 == rd ? _next_reg_T_834[127:64] : _GEN_9053; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9086 = 5'h16 == rd ? _next_reg_T_834[127:64] : _GEN_9054; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9087 = 5'h17 == rd ? _next_reg_T_834[127:64] : _GEN_9055; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9088 = 5'h18 == rd ? _next_reg_T_834[127:64] : _GEN_9056; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9089 = 5'h19 == rd ? _next_reg_T_834[127:64] : _GEN_9057; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9090 = 5'h1a == rd ? _next_reg_T_834[127:64] : _GEN_9058; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9091 = 5'h1b == rd ? _next_reg_T_834[127:64] : _GEN_9059; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9092 = 5'h1c == rd ? _next_reg_T_834[127:64] : _GEN_9060; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9093 = 5'h1d == rd ? _next_reg_T_834[127:64] : _GEN_9061; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9094 = 5'h1e == rd ? _next_reg_T_834[127:64] : _GEN_9062; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9095 = 5'h1f == rd ? _next_reg_T_834[127:64] : _GEN_9063; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:{48,48}]
  wire [63:0] _GEN_9104 = _T_1496 ? _GEN_9065 : _GEN_9033; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9105 = _T_1496 ? _GEN_9066 : _GEN_9034; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9106 = _T_1496 ? _GEN_9067 : _GEN_9035; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9107 = _T_1496 ? _GEN_9068 : _GEN_9036; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9108 = _T_1496 ? _GEN_9069 : _GEN_9037; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9109 = _T_1496 ? _GEN_9070 : _GEN_9038; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9110 = _T_1496 ? _GEN_9071 : _GEN_9039; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9111 = _T_1496 ? _GEN_9072 : _GEN_9040; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9112 = _T_1496 ? _GEN_9073 : _GEN_9041; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9113 = _T_1496 ? _GEN_9074 : _GEN_9042; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9114 = _T_1496 ? _GEN_9075 : _GEN_9043; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9115 = _T_1496 ? _GEN_9076 : _GEN_9044; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9116 = _T_1496 ? _GEN_9077 : _GEN_9045; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9117 = _T_1496 ? _GEN_9078 : _GEN_9046; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9118 = _T_1496 ? _GEN_9079 : _GEN_9047; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9119 = _T_1496 ? _GEN_9080 : _GEN_9048; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9120 = _T_1496 ? _GEN_9081 : _GEN_9049; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9121 = _T_1496 ? _GEN_9082 : _GEN_9050; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9122 = _T_1496 ? _GEN_9083 : _GEN_9051; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9123 = _T_1496 ? _GEN_9084 : _GEN_9052; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9124 = _T_1496 ? _GEN_9085 : _GEN_9053; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9125 = _T_1496 ? _GEN_9086 : _GEN_9054; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9126 = _T_1496 ? _GEN_9087 : _GEN_9055; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9127 = _T_1496 ? _GEN_9088 : _GEN_9056; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9128 = _T_1496 ? _GEN_9089 : _GEN_9057; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9129 = _T_1496 ? _GEN_9090 : _GEN_9058; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9130 = _T_1496 ? _GEN_9091 : _GEN_9059; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9131 = _T_1496 ? _GEN_9092 : _GEN_9060; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9132 = _T_1496 ? _GEN_9093 : _GEN_9061; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9133 = _T_1496 ? _GEN_9094 : _GEN_9062; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [63:0] _GEN_9134 = _T_1496 ? _GEN_9095 : _GEN_9063; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 88:24]
  wire [64:0] _next_reg_T_852 = $signed(_T_325) / $signed(_T_326); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 49:23]
  wire  _next_reg_T_854 = _GEN_910 == 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 51:19]
  wire [63:0] _next_reg_T_858 = 64'h0 - 64'hffffffff80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:22]
  wire  _next_reg_T_862 = _GEN_101 == _next_reg_T_858 & _GEN_910 == 64'hffffffffffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:52]
  wire [63:0] _next_reg_T_866 = _next_reg_T_862 ? _next_reg_T_858 : _next_reg_T_852[63:0]; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _next_reg_T_867 = _next_reg_T_854 ? 64'hffffffffffffffff : _next_reg_T_866; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _GEN_9136 = 5'h1 == rd ? _next_reg_T_867 : _GEN_9104; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9137 = 5'h2 == rd ? _next_reg_T_867 : _GEN_9105; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9138 = 5'h3 == rd ? _next_reg_T_867 : _GEN_9106; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9139 = 5'h4 == rd ? _next_reg_T_867 : _GEN_9107; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9140 = 5'h5 == rd ? _next_reg_T_867 : _GEN_9108; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9141 = 5'h6 == rd ? _next_reg_T_867 : _GEN_9109; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9142 = 5'h7 == rd ? _next_reg_T_867 : _GEN_9110; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9143 = 5'h8 == rd ? _next_reg_T_867 : _GEN_9111; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9144 = 5'h9 == rd ? _next_reg_T_867 : _GEN_9112; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9145 = 5'ha == rd ? _next_reg_T_867 : _GEN_9113; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9146 = 5'hb == rd ? _next_reg_T_867 : _GEN_9114; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9147 = 5'hc == rd ? _next_reg_T_867 : _GEN_9115; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9148 = 5'hd == rd ? _next_reg_T_867 : _GEN_9116; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9149 = 5'he == rd ? _next_reg_T_867 : _GEN_9117; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9150 = 5'hf == rd ? _next_reg_T_867 : _GEN_9118; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9151 = 5'h10 == rd ? _next_reg_T_867 : _GEN_9119; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9152 = 5'h11 == rd ? _next_reg_T_867 : _GEN_9120; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9153 = 5'h12 == rd ? _next_reg_T_867 : _GEN_9121; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9154 = 5'h13 == rd ? _next_reg_T_867 : _GEN_9122; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9155 = 5'h14 == rd ? _next_reg_T_867 : _GEN_9123; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9156 = 5'h15 == rd ? _next_reg_T_867 : _GEN_9124; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9157 = 5'h16 == rd ? _next_reg_T_867 : _GEN_9125; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9158 = 5'h17 == rd ? _next_reg_T_867 : _GEN_9126; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9159 = 5'h18 == rd ? _next_reg_T_867 : _GEN_9127; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9160 = 5'h19 == rd ? _next_reg_T_867 : _GEN_9128; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9161 = 5'h1a == rd ? _next_reg_T_867 : _GEN_9129; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9162 = 5'h1b == rd ? _next_reg_T_867 : _GEN_9130; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9163 = 5'h1c == rd ? _next_reg_T_867 : _GEN_9131; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9164 = 5'h1d == rd ? _next_reg_T_867 : _GEN_9132; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9165 = 5'h1e == rd ? _next_reg_T_867 : _GEN_9133; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9166 = 5'h1f == rd ? _next_reg_T_867 : _GEN_9134; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:{46,46}]
  wire [63:0] _GEN_9175 = _T_1503 ? _GEN_9136 : _GEN_9104; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9176 = _T_1503 ? _GEN_9137 : _GEN_9105; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9177 = _T_1503 ? _GEN_9138 : _GEN_9106; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9178 = _T_1503 ? _GEN_9139 : _GEN_9107; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9179 = _T_1503 ? _GEN_9140 : _GEN_9108; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9180 = _T_1503 ? _GEN_9141 : _GEN_9109; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9181 = _T_1503 ? _GEN_9142 : _GEN_9110; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9182 = _T_1503 ? _GEN_9143 : _GEN_9111; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9183 = _T_1503 ? _GEN_9144 : _GEN_9112; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9184 = _T_1503 ? _GEN_9145 : _GEN_9113; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9185 = _T_1503 ? _GEN_9146 : _GEN_9114; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9186 = _T_1503 ? _GEN_9147 : _GEN_9115; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9187 = _T_1503 ? _GEN_9148 : _GEN_9116; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9188 = _T_1503 ? _GEN_9149 : _GEN_9117; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9189 = _T_1503 ? _GEN_9150 : _GEN_9118; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9190 = _T_1503 ? _GEN_9151 : _GEN_9119; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9191 = _T_1503 ? _GEN_9152 : _GEN_9120; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9192 = _T_1503 ? _GEN_9153 : _GEN_9121; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9193 = _T_1503 ? _GEN_9154 : _GEN_9122; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9194 = _T_1503 ? _GEN_9155 : _GEN_9123; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9195 = _T_1503 ? _GEN_9156 : _GEN_9124; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9196 = _T_1503 ? _GEN_9157 : _GEN_9125; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9197 = _T_1503 ? _GEN_9158 : _GEN_9126; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9198 = _T_1503 ? _GEN_9159 : _GEN_9127; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9199 = _T_1503 ? _GEN_9160 : _GEN_9128; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9200 = _T_1503 ? _GEN_9161 : _GEN_9129; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9201 = _T_1503 ? _GEN_9162 : _GEN_9130; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9202 = _T_1503 ? _GEN_9163 : _GEN_9131; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9203 = _T_1503 ? _GEN_9164 : _GEN_9132; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9204 = _T_1503 ? _GEN_9165 : _GEN_9133; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _GEN_9205 = _T_1503 ? _GEN_9166 : _GEN_9134; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 91:22]
  wire [63:0] _next_reg_T_868 = _GEN_101 / _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 58:15]
  wire [63:0] _next_reg_T_871 = _next_reg_T_854 ? 64'hffffffffffffffff : _next_reg_T_868; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _GEN_9207 = 5'h1 == rd ? _next_reg_T_871 : _GEN_9175; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9208 = 5'h2 == rd ? _next_reg_T_871 : _GEN_9176; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9209 = 5'h3 == rd ? _next_reg_T_871 : _GEN_9177; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9210 = 5'h4 == rd ? _next_reg_T_871 : _GEN_9178; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9211 = 5'h5 == rd ? _next_reg_T_871 : _GEN_9179; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9212 = 5'h6 == rd ? _next_reg_T_871 : _GEN_9180; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9213 = 5'h7 == rd ? _next_reg_T_871 : _GEN_9181; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9214 = 5'h8 == rd ? _next_reg_T_871 : _GEN_9182; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9215 = 5'h9 == rd ? _next_reg_T_871 : _GEN_9183; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9216 = 5'ha == rd ? _next_reg_T_871 : _GEN_9184; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9217 = 5'hb == rd ? _next_reg_T_871 : _GEN_9185; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9218 = 5'hc == rd ? _next_reg_T_871 : _GEN_9186; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9219 = 5'hd == rd ? _next_reg_T_871 : _GEN_9187; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9220 = 5'he == rd ? _next_reg_T_871 : _GEN_9188; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9221 = 5'hf == rd ? _next_reg_T_871 : _GEN_9189; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9222 = 5'h10 == rd ? _next_reg_T_871 : _GEN_9190; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9223 = 5'h11 == rd ? _next_reg_T_871 : _GEN_9191; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9224 = 5'h12 == rd ? _next_reg_T_871 : _GEN_9192; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9225 = 5'h13 == rd ? _next_reg_T_871 : _GEN_9193; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9226 = 5'h14 == rd ? _next_reg_T_871 : _GEN_9194; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9227 = 5'h15 == rd ? _next_reg_T_871 : _GEN_9195; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9228 = 5'h16 == rd ? _next_reg_T_871 : _GEN_9196; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9229 = 5'h17 == rd ? _next_reg_T_871 : _GEN_9197; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9230 = 5'h18 == rd ? _next_reg_T_871 : _GEN_9198; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9231 = 5'h19 == rd ? _next_reg_T_871 : _GEN_9199; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9232 = 5'h1a == rd ? _next_reg_T_871 : _GEN_9200; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9233 = 5'h1b == rd ? _next_reg_T_871 : _GEN_9201; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9234 = 5'h1c == rd ? _next_reg_T_871 : _GEN_9202; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9235 = 5'h1d == rd ? _next_reg_T_871 : _GEN_9203; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9236 = 5'h1e == rd ? _next_reg_T_871 : _GEN_9204; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9237 = 5'h1f == rd ? _next_reg_T_871 : _GEN_9205; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:{46,46}]
  wire [63:0] _GEN_9246 = _T_1510 ? _GEN_9207 : _GEN_9175; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9247 = _T_1510 ? _GEN_9208 : _GEN_9176; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9248 = _T_1510 ? _GEN_9209 : _GEN_9177; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9249 = _T_1510 ? _GEN_9210 : _GEN_9178; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9250 = _T_1510 ? _GEN_9211 : _GEN_9179; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9251 = _T_1510 ? _GEN_9212 : _GEN_9180; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9252 = _T_1510 ? _GEN_9213 : _GEN_9181; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9253 = _T_1510 ? _GEN_9214 : _GEN_9182; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9254 = _T_1510 ? _GEN_9215 : _GEN_9183; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9255 = _T_1510 ? _GEN_9216 : _GEN_9184; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9256 = _T_1510 ? _GEN_9217 : _GEN_9185; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9257 = _T_1510 ? _GEN_9218 : _GEN_9186; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9258 = _T_1510 ? _GEN_9219 : _GEN_9187; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9259 = _T_1510 ? _GEN_9220 : _GEN_9188; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9260 = _T_1510 ? _GEN_9221 : _GEN_9189; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9261 = _T_1510 ? _GEN_9222 : _GEN_9190; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9262 = _T_1510 ? _GEN_9223 : _GEN_9191; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9263 = _T_1510 ? _GEN_9224 : _GEN_9192; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9264 = _T_1510 ? _GEN_9225 : _GEN_9193; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9265 = _T_1510 ? _GEN_9226 : _GEN_9194; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9266 = _T_1510 ? _GEN_9227 : _GEN_9195; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9267 = _T_1510 ? _GEN_9228 : _GEN_9196; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9268 = _T_1510 ? _GEN_9229 : _GEN_9197; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9269 = _T_1510 ? _GEN_9230 : _GEN_9198; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9270 = _T_1510 ? _GEN_9231 : _GEN_9199; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9271 = _T_1510 ? _GEN_9232 : _GEN_9200; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9272 = _T_1510 ? _GEN_9233 : _GEN_9201; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9273 = _T_1510 ? _GEN_9234 : _GEN_9202; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9274 = _T_1510 ? _GEN_9235 : _GEN_9203; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9275 = _T_1510 ? _GEN_9236 : _GEN_9204; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _GEN_9276 = _T_1510 ? _GEN_9237 : _GEN_9205; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 92:22]
  wire [63:0] _next_reg_T_875 = $signed(_T_325) % $signed(_T_326); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 66:42]
  wire [63:0] _next_reg_T_884 = _next_reg_T_862 ? 64'h0 : _next_reg_T_875; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _next_reg_T_885 = _next_reg_T_854 ? _GEN_101 : _next_reg_T_884; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _GEN_9278 = 5'h1 == rd ? _next_reg_T_885 : _GEN_9246; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9279 = 5'h2 == rd ? _next_reg_T_885 : _GEN_9247; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9280 = 5'h3 == rd ? _next_reg_T_885 : _GEN_9248; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9281 = 5'h4 == rd ? _next_reg_T_885 : _GEN_9249; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9282 = 5'h5 == rd ? _next_reg_T_885 : _GEN_9250; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9283 = 5'h6 == rd ? _next_reg_T_885 : _GEN_9251; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9284 = 5'h7 == rd ? _next_reg_T_885 : _GEN_9252; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9285 = 5'h8 == rd ? _next_reg_T_885 : _GEN_9253; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9286 = 5'h9 == rd ? _next_reg_T_885 : _GEN_9254; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9287 = 5'ha == rd ? _next_reg_T_885 : _GEN_9255; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9288 = 5'hb == rd ? _next_reg_T_885 : _GEN_9256; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9289 = 5'hc == rd ? _next_reg_T_885 : _GEN_9257; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9290 = 5'hd == rd ? _next_reg_T_885 : _GEN_9258; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9291 = 5'he == rd ? _next_reg_T_885 : _GEN_9259; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9292 = 5'hf == rd ? _next_reg_T_885 : _GEN_9260; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9293 = 5'h10 == rd ? _next_reg_T_885 : _GEN_9261; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9294 = 5'h11 == rd ? _next_reg_T_885 : _GEN_9262; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9295 = 5'h12 == rd ? _next_reg_T_885 : _GEN_9263; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9296 = 5'h13 == rd ? _next_reg_T_885 : _GEN_9264; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9297 = 5'h14 == rd ? _next_reg_T_885 : _GEN_9265; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9298 = 5'h15 == rd ? _next_reg_T_885 : _GEN_9266; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9299 = 5'h16 == rd ? _next_reg_T_885 : _GEN_9267; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9300 = 5'h17 == rd ? _next_reg_T_885 : _GEN_9268; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9301 = 5'h18 == rd ? _next_reg_T_885 : _GEN_9269; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9302 = 5'h19 == rd ? _next_reg_T_885 : _GEN_9270; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9303 = 5'h1a == rd ? _next_reg_T_885 : _GEN_9271; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9304 = 5'h1b == rd ? _next_reg_T_885 : _GEN_9272; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9305 = 5'h1c == rd ? _next_reg_T_885 : _GEN_9273; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9306 = 5'h1d == rd ? _next_reg_T_885 : _GEN_9274; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9307 = 5'h1e == rd ? _next_reg_T_885 : _GEN_9275; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9308 = 5'h1f == rd ? _next_reg_T_885 : _GEN_9276; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:{46,46}]
  wire [63:0] _GEN_9317 = _T_1517 ? _GEN_9278 : _GEN_9246; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9318 = _T_1517 ? _GEN_9279 : _GEN_9247; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9319 = _T_1517 ? _GEN_9280 : _GEN_9248; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9320 = _T_1517 ? _GEN_9281 : _GEN_9249; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9321 = _T_1517 ? _GEN_9282 : _GEN_9250; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9322 = _T_1517 ? _GEN_9283 : _GEN_9251; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9323 = _T_1517 ? _GEN_9284 : _GEN_9252; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9324 = _T_1517 ? _GEN_9285 : _GEN_9253; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9325 = _T_1517 ? _GEN_9286 : _GEN_9254; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9326 = _T_1517 ? _GEN_9287 : _GEN_9255; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9327 = _T_1517 ? _GEN_9288 : _GEN_9256; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9328 = _T_1517 ? _GEN_9289 : _GEN_9257; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9329 = _T_1517 ? _GEN_9290 : _GEN_9258; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9330 = _T_1517 ? _GEN_9291 : _GEN_9259; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9331 = _T_1517 ? _GEN_9292 : _GEN_9260; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9332 = _T_1517 ? _GEN_9293 : _GEN_9261; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9333 = _T_1517 ? _GEN_9294 : _GEN_9262; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9334 = _T_1517 ? _GEN_9295 : _GEN_9263; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9335 = _T_1517 ? _GEN_9296 : _GEN_9264; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9336 = _T_1517 ? _GEN_9297 : _GEN_9265; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9337 = _T_1517 ? _GEN_9298 : _GEN_9266; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9338 = _T_1517 ? _GEN_9299 : _GEN_9267; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9339 = _T_1517 ? _GEN_9300 : _GEN_9268; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9340 = _T_1517 ? _GEN_9301 : _GEN_9269; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9341 = _T_1517 ? _GEN_9302 : _GEN_9270; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9342 = _T_1517 ? _GEN_9303 : _GEN_9271; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9343 = _T_1517 ? _GEN_9304 : _GEN_9272; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9344 = _T_1517 ? _GEN_9305 : _GEN_9273; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9345 = _T_1517 ? _GEN_9306 : _GEN_9274; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9346 = _T_1517 ? _GEN_9307 : _GEN_9275; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _GEN_9347 = _T_1517 ? _GEN_9308 : _GEN_9276; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 93:22]
  wire [63:0] _next_reg_T_886 = _GEN_101 % _GEN_910; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 75:15]
  wire [63:0] _next_reg_T_888 = _next_reg_T_854 ? _GEN_101 : _next_reg_T_886; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [63:0] _GEN_9349 = 5'h1 == rd ? _next_reg_T_888 : _GEN_9317; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9350 = 5'h2 == rd ? _next_reg_T_888 : _GEN_9318; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9351 = 5'h3 == rd ? _next_reg_T_888 : _GEN_9319; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9352 = 5'h4 == rd ? _next_reg_T_888 : _GEN_9320; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9353 = 5'h5 == rd ? _next_reg_T_888 : _GEN_9321; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9354 = 5'h6 == rd ? _next_reg_T_888 : _GEN_9322; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9355 = 5'h7 == rd ? _next_reg_T_888 : _GEN_9323; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9356 = 5'h8 == rd ? _next_reg_T_888 : _GEN_9324; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9357 = 5'h9 == rd ? _next_reg_T_888 : _GEN_9325; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9358 = 5'ha == rd ? _next_reg_T_888 : _GEN_9326; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9359 = 5'hb == rd ? _next_reg_T_888 : _GEN_9327; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9360 = 5'hc == rd ? _next_reg_T_888 : _GEN_9328; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9361 = 5'hd == rd ? _next_reg_T_888 : _GEN_9329; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9362 = 5'he == rd ? _next_reg_T_888 : _GEN_9330; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9363 = 5'hf == rd ? _next_reg_T_888 : _GEN_9331; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9364 = 5'h10 == rd ? _next_reg_T_888 : _GEN_9332; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9365 = 5'h11 == rd ? _next_reg_T_888 : _GEN_9333; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9366 = 5'h12 == rd ? _next_reg_T_888 : _GEN_9334; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9367 = 5'h13 == rd ? _next_reg_T_888 : _GEN_9335; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9368 = 5'h14 == rd ? _next_reg_T_888 : _GEN_9336; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9369 = 5'h15 == rd ? _next_reg_T_888 : _GEN_9337; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9370 = 5'h16 == rd ? _next_reg_T_888 : _GEN_9338; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9371 = 5'h17 == rd ? _next_reg_T_888 : _GEN_9339; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9372 = 5'h18 == rd ? _next_reg_T_888 : _GEN_9340; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9373 = 5'h19 == rd ? _next_reg_T_888 : _GEN_9341; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9374 = 5'h1a == rd ? _next_reg_T_888 : _GEN_9342; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9375 = 5'h1b == rd ? _next_reg_T_888 : _GEN_9343; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9376 = 5'h1c == rd ? _next_reg_T_888 : _GEN_9344; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9377 = 5'h1d == rd ? _next_reg_T_888 : _GEN_9345; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9378 = 5'h1e == rd ? _next_reg_T_888 : _GEN_9346; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9379 = 5'h1f == rd ? _next_reg_T_888 : _GEN_9347; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:{46,46}]
  wire [63:0] _GEN_9388 = _T_1524 ? _GEN_9349 : _GEN_9317; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9389 = _T_1524 ? _GEN_9350 : _GEN_9318; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9390 = _T_1524 ? _GEN_9351 : _GEN_9319; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9391 = _T_1524 ? _GEN_9352 : _GEN_9320; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9392 = _T_1524 ? _GEN_9353 : _GEN_9321; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9393 = _T_1524 ? _GEN_9354 : _GEN_9322; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9394 = _T_1524 ? _GEN_9355 : _GEN_9323; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9395 = _T_1524 ? _GEN_9356 : _GEN_9324; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9396 = _T_1524 ? _GEN_9357 : _GEN_9325; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9397 = _T_1524 ? _GEN_9358 : _GEN_9326; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9398 = _T_1524 ? _GEN_9359 : _GEN_9327; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9399 = _T_1524 ? _GEN_9360 : _GEN_9328; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9400 = _T_1524 ? _GEN_9361 : _GEN_9329; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9401 = _T_1524 ? _GEN_9362 : _GEN_9330; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9402 = _T_1524 ? _GEN_9363 : _GEN_9331; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9403 = _T_1524 ? _GEN_9364 : _GEN_9332; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9404 = _T_1524 ? _GEN_9365 : _GEN_9333; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9405 = _T_1524 ? _GEN_9366 : _GEN_9334; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9406 = _T_1524 ? _GEN_9367 : _GEN_9335; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9407 = _T_1524 ? _GEN_9368 : _GEN_9336; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9408 = _T_1524 ? _GEN_9369 : _GEN_9337; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9409 = _T_1524 ? _GEN_9370 : _GEN_9338; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9410 = _T_1524 ? _GEN_9371 : _GEN_9339; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9411 = _T_1524 ? _GEN_9372 : _GEN_9340; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9412 = _T_1524 ? _GEN_9373 : _GEN_9341; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9413 = _T_1524 ? _GEN_9374 : _GEN_9342; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9414 = _T_1524 ? _GEN_9375 : _GEN_9343; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9415 = _T_1524 ? _GEN_9376 : _GEN_9344; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9416 = _T_1524 ? _GEN_9377 : _GEN_9345; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9417 = _T_1524 ? _GEN_9378 : _GEN_9346; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _GEN_9418 = _T_1524 ? _GEN_9379 : _GEN_9347; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 94:22]
  wire [63:0] _next_reg_T_891 = _GEN_101[31:0] * _GEN_910[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:78]
  wire  next_reg_signBit_20 = _next_reg_T_891[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_894 = next_reg_signBit_20 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_895 = {_next_reg_T_894,_next_reg_T_891[31:0]}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_9420 = 5'h1 == rd ? _next_reg_T_895 : _GEN_9388; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9421 = 5'h2 == rd ? _next_reg_T_895 : _GEN_9389; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9422 = 5'h3 == rd ? _next_reg_T_895 : _GEN_9390; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9423 = 5'h4 == rd ? _next_reg_T_895 : _GEN_9391; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9424 = 5'h5 == rd ? _next_reg_T_895 : _GEN_9392; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9425 = 5'h6 == rd ? _next_reg_T_895 : _GEN_9393; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9426 = 5'h7 == rd ? _next_reg_T_895 : _GEN_9394; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9427 = 5'h8 == rd ? _next_reg_T_895 : _GEN_9395; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9428 = 5'h9 == rd ? _next_reg_T_895 : _GEN_9396; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9429 = 5'ha == rd ? _next_reg_T_895 : _GEN_9397; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9430 = 5'hb == rd ? _next_reg_T_895 : _GEN_9398; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9431 = 5'hc == rd ? _next_reg_T_895 : _GEN_9399; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9432 = 5'hd == rd ? _next_reg_T_895 : _GEN_9400; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9433 = 5'he == rd ? _next_reg_T_895 : _GEN_9401; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9434 = 5'hf == rd ? _next_reg_T_895 : _GEN_9402; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9435 = 5'h10 == rd ? _next_reg_T_895 : _GEN_9403; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9436 = 5'h11 == rd ? _next_reg_T_895 : _GEN_9404; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9437 = 5'h12 == rd ? _next_reg_T_895 : _GEN_9405; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9438 = 5'h13 == rd ? _next_reg_T_895 : _GEN_9406; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9439 = 5'h14 == rd ? _next_reg_T_895 : _GEN_9407; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9440 = 5'h15 == rd ? _next_reg_T_895 : _GEN_9408; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9441 = 5'h16 == rd ? _next_reg_T_895 : _GEN_9409; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9442 = 5'h17 == rd ? _next_reg_T_895 : _GEN_9410; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9443 = 5'h18 == rd ? _next_reg_T_895 : _GEN_9411; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9444 = 5'h19 == rd ? _next_reg_T_895 : _GEN_9412; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9445 = 5'h1a == rd ? _next_reg_T_895 : _GEN_9413; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9446 = 5'h1b == rd ? _next_reg_T_895 : _GEN_9414; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9447 = 5'h1c == rd ? _next_reg_T_895 : _GEN_9415; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9448 = 5'h1d == rd ? _next_reg_T_895 : _GEN_9416; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9449 = 5'h1e == rd ? _next_reg_T_895 : _GEN_9417; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9450 = 5'h1f == rd ? _next_reg_T_895 : _GEN_9418; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:{46,46}]
  wire [63:0] _GEN_9459 = _T_1531 ? _GEN_9420 : _GEN_9388; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9460 = _T_1531 ? _GEN_9421 : _GEN_9389; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9461 = _T_1531 ? _GEN_9422 : _GEN_9390; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9462 = _T_1531 ? _GEN_9423 : _GEN_9391; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9463 = _T_1531 ? _GEN_9424 : _GEN_9392; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9464 = _T_1531 ? _GEN_9425 : _GEN_9393; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9465 = _T_1531 ? _GEN_9426 : _GEN_9394; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9466 = _T_1531 ? _GEN_9427 : _GEN_9395; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9467 = _T_1531 ? _GEN_9428 : _GEN_9396; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9468 = _T_1531 ? _GEN_9429 : _GEN_9397; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9469 = _T_1531 ? _GEN_9430 : _GEN_9398; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9470 = _T_1531 ? _GEN_9431 : _GEN_9399; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9471 = _T_1531 ? _GEN_9432 : _GEN_9400; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9472 = _T_1531 ? _GEN_9433 : _GEN_9401; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9473 = _T_1531 ? _GEN_9434 : _GEN_9402; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9474 = _T_1531 ? _GEN_9435 : _GEN_9403; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9475 = _T_1531 ? _GEN_9436 : _GEN_9404; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9476 = _T_1531 ? _GEN_9437 : _GEN_9405; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9477 = _T_1531 ? _GEN_9438 : _GEN_9406; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9478 = _T_1531 ? _GEN_9439 : _GEN_9407; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9479 = _T_1531 ? _GEN_9440 : _GEN_9408; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9480 = _T_1531 ? _GEN_9441 : _GEN_9409; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9481 = _T_1531 ? _GEN_9442 : _GEN_9410; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9482 = _T_1531 ? _GEN_9443 : _GEN_9411; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9483 = _T_1531 ? _GEN_9444 : _GEN_9412; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9484 = _T_1531 ? _GEN_9445 : _GEN_9413; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9485 = _T_1531 ? _GEN_9446 : _GEN_9414; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9486 = _T_1531 ? _GEN_9447 : _GEN_9415; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9487 = _T_1531 ? _GEN_9448 : _GEN_9416; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9488 = _T_1531 ? _GEN_9449 : _GEN_9417; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [63:0] _GEN_9489 = _T_1531 ? _GEN_9450 : _GEN_9418; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 102:22]
  wire [31:0] _next_reg_T_899 = _GEN_910[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 49:34]
  wire [32:0] _next_reg_T_900 = $signed(_next_reg_T_370) / $signed(_next_reg_T_899); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 49:23]
  wire  _next_reg_T_902 = _GEN_910[31:0] == 32'h0; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 51:19]
  wire [31:0] _next_reg_T_906 = 32'h0 - 32'h80000000; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:22]
  wire  _next_reg_T_910 = _GEN_101[31:0] == _next_reg_T_906 & _GEN_910[31:0] == 32'hffffffff; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 52:52]
  wire [31:0] _next_reg_T_914 = _next_reg_T_910 ? _next_reg_T_906 : _next_reg_T_900[31:0]; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _next_reg_T_915 = _next_reg_T_902 ? 32'hffffffff : _next_reg_T_914; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  next_reg_signBit_21 = _next_reg_T_915[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_917 = next_reg_signBit_21 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_918 = {_next_reg_T_917,_next_reg_T_915}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_9491 = 5'h1 == rd ? _next_reg_T_918 : _GEN_9459; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9492 = 5'h2 == rd ? _next_reg_T_918 : _GEN_9460; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9493 = 5'h3 == rd ? _next_reg_T_918 : _GEN_9461; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9494 = 5'h4 == rd ? _next_reg_T_918 : _GEN_9462; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9495 = 5'h5 == rd ? _next_reg_T_918 : _GEN_9463; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9496 = 5'h6 == rd ? _next_reg_T_918 : _GEN_9464; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9497 = 5'h7 == rd ? _next_reg_T_918 : _GEN_9465; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9498 = 5'h8 == rd ? _next_reg_T_918 : _GEN_9466; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9499 = 5'h9 == rd ? _next_reg_T_918 : _GEN_9467; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9500 = 5'ha == rd ? _next_reg_T_918 : _GEN_9468; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9501 = 5'hb == rd ? _next_reg_T_918 : _GEN_9469; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9502 = 5'hc == rd ? _next_reg_T_918 : _GEN_9470; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9503 = 5'hd == rd ? _next_reg_T_918 : _GEN_9471; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9504 = 5'he == rd ? _next_reg_T_918 : _GEN_9472; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9505 = 5'hf == rd ? _next_reg_T_918 : _GEN_9473; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9506 = 5'h10 == rd ? _next_reg_T_918 : _GEN_9474; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9507 = 5'h11 == rd ? _next_reg_T_918 : _GEN_9475; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9508 = 5'h12 == rd ? _next_reg_T_918 : _GEN_9476; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9509 = 5'h13 == rd ? _next_reg_T_918 : _GEN_9477; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9510 = 5'h14 == rd ? _next_reg_T_918 : _GEN_9478; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9511 = 5'h15 == rd ? _next_reg_T_918 : _GEN_9479; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9512 = 5'h16 == rd ? _next_reg_T_918 : _GEN_9480; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9513 = 5'h17 == rd ? _next_reg_T_918 : _GEN_9481; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9514 = 5'h18 == rd ? _next_reg_T_918 : _GEN_9482; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9515 = 5'h19 == rd ? _next_reg_T_918 : _GEN_9483; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9516 = 5'h1a == rd ? _next_reg_T_918 : _GEN_9484; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9517 = 5'h1b == rd ? _next_reg_T_918 : _GEN_9485; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9518 = 5'h1c == rd ? _next_reg_T_918 : _GEN_9486; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9519 = 5'h1d == rd ? _next_reg_T_918 : _GEN_9487; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9520 = 5'h1e == rd ? _next_reg_T_918 : _GEN_9488; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9521 = 5'h1f == rd ? _next_reg_T_918 : _GEN_9489; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:{47,47}]
  wire [63:0] _GEN_9530 = _T_1538 ? _GEN_9491 : _GEN_9459; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9531 = _T_1538 ? _GEN_9492 : _GEN_9460; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9532 = _T_1538 ? _GEN_9493 : _GEN_9461; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9533 = _T_1538 ? _GEN_9494 : _GEN_9462; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9534 = _T_1538 ? _GEN_9495 : _GEN_9463; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9535 = _T_1538 ? _GEN_9496 : _GEN_9464; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9536 = _T_1538 ? _GEN_9497 : _GEN_9465; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9537 = _T_1538 ? _GEN_9498 : _GEN_9466; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9538 = _T_1538 ? _GEN_9499 : _GEN_9467; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9539 = _T_1538 ? _GEN_9500 : _GEN_9468; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9540 = _T_1538 ? _GEN_9501 : _GEN_9469; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9541 = _T_1538 ? _GEN_9502 : _GEN_9470; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9542 = _T_1538 ? _GEN_9503 : _GEN_9471; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9543 = _T_1538 ? _GEN_9504 : _GEN_9472; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9544 = _T_1538 ? _GEN_9505 : _GEN_9473; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9545 = _T_1538 ? _GEN_9506 : _GEN_9474; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9546 = _T_1538 ? _GEN_9507 : _GEN_9475; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9547 = _T_1538 ? _GEN_9508 : _GEN_9476; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9548 = _T_1538 ? _GEN_9509 : _GEN_9477; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9549 = _T_1538 ? _GEN_9510 : _GEN_9478; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9550 = _T_1538 ? _GEN_9511 : _GEN_9479; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9551 = _T_1538 ? _GEN_9512 : _GEN_9480; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9552 = _T_1538 ? _GEN_9513 : _GEN_9481; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9553 = _T_1538 ? _GEN_9514 : _GEN_9482; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9554 = _T_1538 ? _GEN_9515 : _GEN_9483; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9555 = _T_1538 ? _GEN_9516 : _GEN_9484; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9556 = _T_1538 ? _GEN_9517 : _GEN_9485; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9557 = _T_1538 ? _GEN_9518 : _GEN_9486; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9558 = _T_1538 ? _GEN_9519 : _GEN_9487; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9559 = _T_1538 ? _GEN_9520 : _GEN_9488; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [63:0] _GEN_9560 = _T_1538 ? _GEN_9521 : _GEN_9489; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 105:23]
  wire [31:0] _next_reg_T_921 = _GEN_101[31:0] / _GEN_910[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 58:15]
  wire [31:0] _next_reg_T_924 = _next_reg_T_902 ? 32'hffffffff : _next_reg_T_921; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  next_reg_signBit_22 = _next_reg_T_924[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_926 = next_reg_signBit_22 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_927 = {_next_reg_T_926,_next_reg_T_924}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_9562 = 5'h1 == rd ? _next_reg_T_927 : _GEN_9530; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9563 = 5'h2 == rd ? _next_reg_T_927 : _GEN_9531; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9564 = 5'h3 == rd ? _next_reg_T_927 : _GEN_9532; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9565 = 5'h4 == rd ? _next_reg_T_927 : _GEN_9533; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9566 = 5'h5 == rd ? _next_reg_T_927 : _GEN_9534; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9567 = 5'h6 == rd ? _next_reg_T_927 : _GEN_9535; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9568 = 5'h7 == rd ? _next_reg_T_927 : _GEN_9536; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9569 = 5'h8 == rd ? _next_reg_T_927 : _GEN_9537; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9570 = 5'h9 == rd ? _next_reg_T_927 : _GEN_9538; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9571 = 5'ha == rd ? _next_reg_T_927 : _GEN_9539; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9572 = 5'hb == rd ? _next_reg_T_927 : _GEN_9540; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9573 = 5'hc == rd ? _next_reg_T_927 : _GEN_9541; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9574 = 5'hd == rd ? _next_reg_T_927 : _GEN_9542; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9575 = 5'he == rd ? _next_reg_T_927 : _GEN_9543; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9576 = 5'hf == rd ? _next_reg_T_927 : _GEN_9544; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9577 = 5'h10 == rd ? _next_reg_T_927 : _GEN_9545; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9578 = 5'h11 == rd ? _next_reg_T_927 : _GEN_9546; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9579 = 5'h12 == rd ? _next_reg_T_927 : _GEN_9547; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9580 = 5'h13 == rd ? _next_reg_T_927 : _GEN_9548; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9581 = 5'h14 == rd ? _next_reg_T_927 : _GEN_9549; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9582 = 5'h15 == rd ? _next_reg_T_927 : _GEN_9550; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9583 = 5'h16 == rd ? _next_reg_T_927 : _GEN_9551; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9584 = 5'h17 == rd ? _next_reg_T_927 : _GEN_9552; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9585 = 5'h18 == rd ? _next_reg_T_927 : _GEN_9553; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9586 = 5'h19 == rd ? _next_reg_T_927 : _GEN_9554; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9587 = 5'h1a == rd ? _next_reg_T_927 : _GEN_9555; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9588 = 5'h1b == rd ? _next_reg_T_927 : _GEN_9556; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9589 = 5'h1c == rd ? _next_reg_T_927 : _GEN_9557; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9590 = 5'h1d == rd ? _next_reg_T_927 : _GEN_9558; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9591 = 5'h1e == rd ? _next_reg_T_927 : _GEN_9559; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9592 = 5'h1f == rd ? _next_reg_T_927 : _GEN_9560; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:{47,47}]
  wire [63:0] _GEN_9601 = _T_1545 ? _GEN_9562 : _GEN_9530; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9602 = _T_1545 ? _GEN_9563 : _GEN_9531; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9603 = _T_1545 ? _GEN_9564 : _GEN_9532; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9604 = _T_1545 ? _GEN_9565 : _GEN_9533; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9605 = _T_1545 ? _GEN_9566 : _GEN_9534; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9606 = _T_1545 ? _GEN_9567 : _GEN_9535; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9607 = _T_1545 ? _GEN_9568 : _GEN_9536; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9608 = _T_1545 ? _GEN_9569 : _GEN_9537; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9609 = _T_1545 ? _GEN_9570 : _GEN_9538; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9610 = _T_1545 ? _GEN_9571 : _GEN_9539; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9611 = _T_1545 ? _GEN_9572 : _GEN_9540; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9612 = _T_1545 ? _GEN_9573 : _GEN_9541; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9613 = _T_1545 ? _GEN_9574 : _GEN_9542; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9614 = _T_1545 ? _GEN_9575 : _GEN_9543; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9615 = _T_1545 ? _GEN_9576 : _GEN_9544; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9616 = _T_1545 ? _GEN_9577 : _GEN_9545; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9617 = _T_1545 ? _GEN_9578 : _GEN_9546; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9618 = _T_1545 ? _GEN_9579 : _GEN_9547; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9619 = _T_1545 ? _GEN_9580 : _GEN_9548; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9620 = _T_1545 ? _GEN_9581 : _GEN_9549; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9621 = _T_1545 ? _GEN_9582 : _GEN_9550; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9622 = _T_1545 ? _GEN_9583 : _GEN_9551; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9623 = _T_1545 ? _GEN_9584 : _GEN_9552; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9624 = _T_1545 ? _GEN_9585 : _GEN_9553; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9625 = _T_1545 ? _GEN_9586 : _GEN_9554; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9626 = _T_1545 ? _GEN_9587 : _GEN_9555; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9627 = _T_1545 ? _GEN_9588 : _GEN_9556; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9628 = _T_1545 ? _GEN_9589 : _GEN_9557; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9629 = _T_1545 ? _GEN_9590 : _GEN_9558; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9630 = _T_1545 ? _GEN_9591 : _GEN_9559; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [63:0] _GEN_9631 = _T_1545 ? _GEN_9592 : _GEN_9560; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 106:23]
  wire [31:0] _next_reg_T_933 = $signed(_next_reg_T_370) % $signed(_next_reg_T_899); // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 66:42]
  wire [31:0] _next_reg_T_942 = _next_reg_T_910 ? 32'h0 : _next_reg_T_933; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire [31:0] _next_reg_T_943 = _next_reg_T_902 ? _GEN_101[31:0] : _next_reg_T_942; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  next_reg_signBit_23 = _next_reg_T_943[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_945 = next_reg_signBit_23 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_946 = {_next_reg_T_945,_next_reg_T_943}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_9633 = 5'h1 == rd ? _next_reg_T_946 : _GEN_9601; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9634 = 5'h2 == rd ? _next_reg_T_946 : _GEN_9602; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9635 = 5'h3 == rd ? _next_reg_T_946 : _GEN_9603; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9636 = 5'h4 == rd ? _next_reg_T_946 : _GEN_9604; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9637 = 5'h5 == rd ? _next_reg_T_946 : _GEN_9605; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9638 = 5'h6 == rd ? _next_reg_T_946 : _GEN_9606; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9639 = 5'h7 == rd ? _next_reg_T_946 : _GEN_9607; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9640 = 5'h8 == rd ? _next_reg_T_946 : _GEN_9608; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9641 = 5'h9 == rd ? _next_reg_T_946 : _GEN_9609; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9642 = 5'ha == rd ? _next_reg_T_946 : _GEN_9610; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9643 = 5'hb == rd ? _next_reg_T_946 : _GEN_9611; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9644 = 5'hc == rd ? _next_reg_T_946 : _GEN_9612; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9645 = 5'hd == rd ? _next_reg_T_946 : _GEN_9613; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9646 = 5'he == rd ? _next_reg_T_946 : _GEN_9614; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9647 = 5'hf == rd ? _next_reg_T_946 : _GEN_9615; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9648 = 5'h10 == rd ? _next_reg_T_946 : _GEN_9616; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9649 = 5'h11 == rd ? _next_reg_T_946 : _GEN_9617; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9650 = 5'h12 == rd ? _next_reg_T_946 : _GEN_9618; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9651 = 5'h13 == rd ? _next_reg_T_946 : _GEN_9619; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9652 = 5'h14 == rd ? _next_reg_T_946 : _GEN_9620; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9653 = 5'h15 == rd ? _next_reg_T_946 : _GEN_9621; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9654 = 5'h16 == rd ? _next_reg_T_946 : _GEN_9622; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9655 = 5'h17 == rd ? _next_reg_T_946 : _GEN_9623; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9656 = 5'h18 == rd ? _next_reg_T_946 : _GEN_9624; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9657 = 5'h19 == rd ? _next_reg_T_946 : _GEN_9625; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9658 = 5'h1a == rd ? _next_reg_T_946 : _GEN_9626; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9659 = 5'h1b == rd ? _next_reg_T_946 : _GEN_9627; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9660 = 5'h1c == rd ? _next_reg_T_946 : _GEN_9628; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9661 = 5'h1d == rd ? _next_reg_T_946 : _GEN_9629; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9662 = 5'h1e == rd ? _next_reg_T_946 : _GEN_9630; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9663 = 5'h1f == rd ? _next_reg_T_946 : _GEN_9631; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:{47,47}]
  wire [63:0] _GEN_9672 = _T_1552 ? _GEN_9633 : _GEN_9601; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9673 = _T_1552 ? _GEN_9634 : _GEN_9602; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9674 = _T_1552 ? _GEN_9635 : _GEN_9603; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9675 = _T_1552 ? _GEN_9636 : _GEN_9604; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9676 = _T_1552 ? _GEN_9637 : _GEN_9605; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9677 = _T_1552 ? _GEN_9638 : _GEN_9606; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9678 = _T_1552 ? _GEN_9639 : _GEN_9607; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9679 = _T_1552 ? _GEN_9640 : _GEN_9608; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9680 = _T_1552 ? _GEN_9641 : _GEN_9609; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9681 = _T_1552 ? _GEN_9642 : _GEN_9610; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9682 = _T_1552 ? _GEN_9643 : _GEN_9611; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9683 = _T_1552 ? _GEN_9644 : _GEN_9612; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9684 = _T_1552 ? _GEN_9645 : _GEN_9613; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9685 = _T_1552 ? _GEN_9646 : _GEN_9614; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9686 = _T_1552 ? _GEN_9647 : _GEN_9615; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9687 = _T_1552 ? _GEN_9648 : _GEN_9616; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9688 = _T_1552 ? _GEN_9649 : _GEN_9617; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9689 = _T_1552 ? _GEN_9650 : _GEN_9618; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9690 = _T_1552 ? _GEN_9651 : _GEN_9619; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9691 = _T_1552 ? _GEN_9652 : _GEN_9620; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9692 = _T_1552 ? _GEN_9653 : _GEN_9621; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9693 = _T_1552 ? _GEN_9654 : _GEN_9622; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9694 = _T_1552 ? _GEN_9655 : _GEN_9623; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9695 = _T_1552 ? _GEN_9656 : _GEN_9624; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9696 = _T_1552 ? _GEN_9657 : _GEN_9625; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9697 = _T_1552 ? _GEN_9658 : _GEN_9626; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9698 = _T_1552 ? _GEN_9659 : _GEN_9627; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9699 = _T_1552 ? _GEN_9660 : _GEN_9628; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9700 = _T_1552 ? _GEN_9661 : _GEN_9629; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9701 = _T_1552 ? _GEN_9662 : _GEN_9630; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [63:0] _GEN_9702 = _T_1552 ? _GEN_9663 : _GEN_9631; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 107:23]
  wire [31:0] _next_reg_T_949 = _GEN_101[31:0] % _GEN_910[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 75:15]
  wire [31:0] _next_reg_T_951 = _next_reg_T_902 ? _GEN_101[31:0] : _next_reg_T_949; // @[src/main/scala/chisel3/util/Mux.scala 141:16]
  wire  next_reg_signBit_24 = _next_reg_T_951[31]; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 9:20]
  wire [31:0] _next_reg_T_953 = next_reg_signBit_24 ? 32'hffffffff : 32'h0; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:15]
  wire [63:0] _next_reg_T_954 = {_next_reg_T_953,_next_reg_T_951}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 13:10]
  wire [63:0] _GEN_9704 = 5'h1 == rd ? _next_reg_T_954 : _GEN_9672; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9705 = 5'h2 == rd ? _next_reg_T_954 : _GEN_9673; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9706 = 5'h3 == rd ? _next_reg_T_954 : _GEN_9674; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9707 = 5'h4 == rd ? _next_reg_T_954 : _GEN_9675; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9708 = 5'h5 == rd ? _next_reg_T_954 : _GEN_9676; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9709 = 5'h6 == rd ? _next_reg_T_954 : _GEN_9677; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9710 = 5'h7 == rd ? _next_reg_T_954 : _GEN_9678; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9711 = 5'h8 == rd ? _next_reg_T_954 : _GEN_9679; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9712 = 5'h9 == rd ? _next_reg_T_954 : _GEN_9680; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9713 = 5'ha == rd ? _next_reg_T_954 : _GEN_9681; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9714 = 5'hb == rd ? _next_reg_T_954 : _GEN_9682; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9715 = 5'hc == rd ? _next_reg_T_954 : _GEN_9683; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9716 = 5'hd == rd ? _next_reg_T_954 : _GEN_9684; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9717 = 5'he == rd ? _next_reg_T_954 : _GEN_9685; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9718 = 5'hf == rd ? _next_reg_T_954 : _GEN_9686; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9719 = 5'h10 == rd ? _next_reg_T_954 : _GEN_9687; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9720 = 5'h11 == rd ? _next_reg_T_954 : _GEN_9688; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9721 = 5'h12 == rd ? _next_reg_T_954 : _GEN_9689; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9722 = 5'h13 == rd ? _next_reg_T_954 : _GEN_9690; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9723 = 5'h14 == rd ? _next_reg_T_954 : _GEN_9691; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9724 = 5'h15 == rd ? _next_reg_T_954 : _GEN_9692; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9725 = 5'h16 == rd ? _next_reg_T_954 : _GEN_9693; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9726 = 5'h17 == rd ? _next_reg_T_954 : _GEN_9694; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9727 = 5'h18 == rd ? _next_reg_T_954 : _GEN_9695; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9728 = 5'h19 == rd ? _next_reg_T_954 : _GEN_9696; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9729 = 5'h1a == rd ? _next_reg_T_954 : _GEN_9697; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9730 = 5'h1b == rd ? _next_reg_T_954 : _GEN_9698; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9731 = 5'h1c == rd ? _next_reg_T_954 : _GEN_9699; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9732 = 5'h1d == rd ? _next_reg_T_954 : _GEN_9700; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9733 = 5'h1e == rd ? _next_reg_T_954 : _GEN_9701; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9734 = 5'h1f == rd ? _next_reg_T_954 : _GEN_9702; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:{47,47}]
  wire [63:0] _GEN_9743 = _T_1559 ? _GEN_9704 : _GEN_9672; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9744 = _T_1559 ? _GEN_9705 : _GEN_9673; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9745 = _T_1559 ? _GEN_9706 : _GEN_9674; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9746 = _T_1559 ? _GEN_9707 : _GEN_9675; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9747 = _T_1559 ? _GEN_9708 : _GEN_9676; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9748 = _T_1559 ? _GEN_9709 : _GEN_9677; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9749 = _T_1559 ? _GEN_9710 : _GEN_9678; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9750 = _T_1559 ? _GEN_9711 : _GEN_9679; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9751 = _T_1559 ? _GEN_9712 : _GEN_9680; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9752 = _T_1559 ? _GEN_9713 : _GEN_9681; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9753 = _T_1559 ? _GEN_9714 : _GEN_9682; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9754 = _T_1559 ? _GEN_9715 : _GEN_9683; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9755 = _T_1559 ? _GEN_9716 : _GEN_9684; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9756 = _T_1559 ? _GEN_9717 : _GEN_9685; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9757 = _T_1559 ? _GEN_9718 : _GEN_9686; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9758 = _T_1559 ? _GEN_9719 : _GEN_9687; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9759 = _T_1559 ? _GEN_9720 : _GEN_9688; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9760 = _T_1559 ? _GEN_9721 : _GEN_9689; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9761 = _T_1559 ? _GEN_9722 : _GEN_9690; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9762 = _T_1559 ? _GEN_9723 : _GEN_9691; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9763 = _T_1559 ? _GEN_9724 : _GEN_9692; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9764 = _T_1559 ? _GEN_9725 : _GEN_9693; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9765 = _T_1559 ? _GEN_9726 : _GEN_9694; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9766 = _T_1559 ? _GEN_9727 : _GEN_9695; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9767 = _T_1559 ? _GEN_9728 : _GEN_9696; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9768 = _T_1559 ? _GEN_9729 : _GEN_9697; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9769 = _T_1559 ? _GEN_9730 : _GEN_9698; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9770 = _T_1559 ? _GEN_9731 : _GEN_9699; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9771 = _T_1559 ? _GEN_9732 : _GEN_9700; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9772 = _T_1559 ? _GEN_9733 : _GEN_9701; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [63:0] _GEN_9773 = _T_1559 ? _GEN_9734 : _GEN_9702; // @[src/main/scala/rvspeccore/core/spec/instset/MExtension.scala 108:23]
  wire [1:0] _next_internal_privilegeMode_T = {1'h0,io_now_csr_mstatus[8]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 125:41]
  wire  mstatusNew_sie = illegalSret | illegalSModeSret ? io_now_csr_mstatus[1] : io_now_csr_mstatus[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 124:35]
  wire  mstatusNew_spie = illegalSret | illegalSModeSret ? io_now_csr_mstatus[5] : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 126:35]
  wire [5:0] next_csr_mstatus_lo_lo = {mstatusNew_spie,io_now_csr_mstatus[4],io_now_csr_mstatus[3],io_now_csr_mstatus[2]
    ,mstatusNew_sie,io_now_csr_mstatus[0]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  mstatusNew_spp = (illegalSret | illegalSModeSret) & io_now_csr_mstatus[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 127:35]
  wire [16:0] next_csr_mstatus_lo = {io_now_csr_mstatus[16:15],io_now_csr_mstatus[14:13],next_reg_mstatusStruct_10_mpp,
    io_now_csr_mstatus[10:9],mstatusNew_spp,io_now_csr_mstatus[7],io_now_csr_mstatus[6],next_csr_mstatus_lo_lo}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  mstatusNew_mprv = (illegalSret | illegalSModeSret) & next_reg_mstatusStruct_10_mprv; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 112:30 120:43 128:35]
  wire [5:0] next_csr_mstatus_hi_lo = {mstatusOld_tsr,io_now_csr_mstatus[21],io_now_csr_mstatus[20],
    next_reg_mstatus_mxr_10,io_now_csr_mstatus[18],mstatusNew_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire [63:0] _next_csr_mstatus_T = {io_now_csr_mstatus[63],io_now_csr_mstatus[62:38],io_now_csr_mstatus[37],
    io_now_csr_mstatus[36],io_now_csr_mstatus[35:34],io_now_csr_mstatus[33:32],io_now_csr_mstatus[31:23],
    next_csr_mstatus_hi_lo,next_csr_mstatus_lo}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 129:49]
  wire  _GEN_9775 = illegalSret | illegalSModeSret | _GEN_8506; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_9793 = _T_1566 ? _GEN_9775 : _GEN_8506; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire  _GEN_9805 = io_now_internal_privilegeMode == 2'h3 ? _GEN_9793 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 88:48 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_9819 = _T_1573 ? _GEN_9805 : _GEN_9793; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire  _GEN_9835 = isIllegalAccess_5 | ~has_15 | _GEN_9819; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_9929 = has_15 ? _GEN_9835 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_9973 = _T_1793 ? _GEN_9929 : _GEN_9835; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire  _GEN_9983 = _T_1592 ? _GEN_9973 : _GEN_9819; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire  _GEN_10027 = isIllegalAccess_4 | ~has_15 | _GEN_9983; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_10097 = has_15 ? _GEN_10027 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_10109 = _T_1794 ? _GEN_10097 : _GEN_10027; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire  _GEN_10153 = _T_1751 ? _GEN_10109 : _GEN_10027; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire  _GEN_10163 = _T_1625 ? _GEN_10153 : _GEN_9983; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire  _GEN_10207 = isIllegalAccess_5 | ~has_15 | _GEN_10163; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_10277 = has_15 ? _GEN_10207 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_10289 = _T_1794 ? _GEN_10277 : _GEN_10207; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire  _GEN_10333 = _T_1793 ? _GEN_10289 : _GEN_10207; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire  _GEN_10343 = _T_1667 ? _GEN_10333 : _GEN_10163; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire  _GEN_10387 = isIllegalAccess_5 | ~has_15 | _GEN_10343; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_10481 = has_15 ? _GEN_10387 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_10525 = _T_1793 ? _GEN_10481 : _GEN_10387; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire  _GEN_10535 = _T_1709 ? _GEN_10525 : _GEN_10343; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire  _GEN_10579 = isIllegalAccess_4 | ~has_15 | _GEN_10535; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_10649 = has_15 ? _GEN_10579 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_10661 = _T_1794 ? _GEN_10649 : _GEN_10579; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire  _GEN_10705 = ~isIllegalWrite_4 ? _GEN_10661 : _GEN_10579; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire  _GEN_10715 = _T_1743 ? _GEN_10705 : _GEN_10535; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire  _GEN_10759 = isIllegalAccess_5 | ~has_15 | _GEN_10715; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 76:35 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_10829 = has_15 ? _GEN_10759 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 145:33]
  wire  _GEN_10841 = rs1 != 5'h0 ? _GEN_10829 : _GEN_10759; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire  _GEN_10885 = ~isIllegalWrite_5 ? _GEN_10841 : _GEN_10759; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire  _GEN_10895 = _T_1786 ? _GEN_10885 : _GEN_10715; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire  _GEN_10940 = illegalInstruction | _GEN_10895; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 133:30 145:33]
  wire  raiseExceptionIntr = io_valid & _GEN_10940; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 118:36]
  wire [63:0] _delegS_T = io_now_csr_medeleg >> exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 155:24]
  wire  delegS = _delegS_T[0] & _vmEnable_T_4; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 155:39]
  wire  _T_1829 = 8'h20 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire  _T_1846 = 8'h40 == io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire [63:0] _GEN_10968 = 8'h40 == io_now_csr_MXLEN ? io_now_pc : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 254:35]
  wire [63:0] _GEN_10978 = 8'h20 == io_now_csr_MXLEN ? io_now_pc : _GEN_10968; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 254:35]
  wire [63:0] _GEN_11033 = delegS ? _GEN_10978 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [63:0] _GEN_11050 = raiseExceptionIntr ? _GEN_11033 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [1:0] _GEN_9777 = illegalSret | illegalSModeSret ? io_now_internal_privilegeMode : _next_internal_privilegeMode_T
    ; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 125:35]
  wire [63:0] _GEN_9781 = illegalSret | illegalSModeSret ? io_now_csr_mstatus : _next_csr_mstatus_T; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 129:35]
  wire  _GEN_9783 = illegalSret | illegalSModeSret ? _GEN_6337 : 1'h1; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 132:25]
  wire [63:0] _GEN_9784 = illegalSret | illegalSModeSret ? _GEN_6338 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 120:43 133:25]
  wire [1:0] _GEN_9794 = _T_1566 ? _GEN_9777 : io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [63:0] _GEN_9795 = _T_1566 ? _GEN_9781 : io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire  _GEN_9797 = _T_1566 ? _GEN_9783 : _GEN_6337; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [63:0] _GEN_9798 = _T_1566 ? _GEN_9784 : _GEN_6338; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 50:22]
  wire [5:0] next_csr_mstatus_lo_lo_1 = {io_now_csr_mstatus[5],io_now_csr_mstatus[4],io_now_csr_mstatus[7],
    io_now_csr_mstatus[2],io_now_csr_mstatus[1],io_now_csr_mstatus[0]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [16:0] next_csr_mstatus_lo_1 = {io_now_csr_mstatus[16:15],io_now_csr_mstatus[14:13],2'h0,io_now_csr_mstatus[10:9]
    ,io_now_csr_mstatus[8],1'h1,io_now_csr_mstatus[6],next_csr_mstatus_lo_lo_1}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [5:0] next_csr_mstatus_hi_lo_1 = {mstatusOld_tsr,io_now_csr_mstatus[21],io_now_csr_mstatus[20],
    next_reg_mstatus_mxr_10,io_now_csr_mstatus[18],next_reg_mstatusStruct_10_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [63:0] _next_csr_mstatus_T_1 = {io_now_csr_mstatus[63],io_now_csr_mstatus[62:38],io_now_csr_mstatus[37],
    io_now_csr_mstatus[36],io_now_csr_mstatus[35:34],io_now_csr_mstatus[33:32],io_now_csr_mstatus[31:23],
    next_csr_mstatus_hi_lo_1,next_csr_mstatus_lo_1}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:38]
  wire [31:0] _rData_T_41 = 32'hfffffffc & io_now_csr_mepc[31:0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:63]
  wire [63:0] _nowCSR_T_82 = _has_T_405 ? io_now_csr_misa : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [63:0] _nowCSR_T_84 = _has_T_407 ? io_now_csr_mvendorid : _nowCSR_T_82; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [63:0] _nowCSR_T_86 = _has_T_409 ? io_now_csr_marchid : _nowCSR_T_84; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [63:0] _nowCSR_T_88 = _has_T_411 ? io_now_csr_mimpid : _nowCSR_T_86; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [63:0] _nowCSR_T_90 = _has_T_413 ? io_now_csr_mhartid : _nowCSR_T_88; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [63:0] _nowCSR_T_92 = _has_T_415 ? io_now_csr_mstatus : _nowCSR_T_90; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [63:0] _nowCSR_T_94 = _has_T_417 ? io_now_csr_mscratch : _nowCSR_T_92; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [63:0] _nowCSR_T_96 = _has_T_419 ? io_now_csr_mtvec : _nowCSR_T_94; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [63:0] _nowCSR_T_98 = _has_T_421 ? io_now_csr_mcounteren : _nowCSR_T_96; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [63:0] _nowCSR_T_100 = _has_T_423 ? io_now_csr_mip : _nowCSR_T_98; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [63:0] _nowCSR_T_102 = _has_T_425 ? io_now_csr_mie : _nowCSR_T_100; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [63:0] _nowCSR_T_104 = _has_T_427 ? io_now_csr_mepc : _nowCSR_T_102; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [63:0] _nowCSR_T_106 = _has_T_429 ? io_now_csr_mcause : _nowCSR_T_104; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [63:0] nowCSR_3 = _has_T_431 ? io_now_csr_mtval : _nowCSR_T_106; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 24:44]
  wire [63:0] _rmask_T_138 = _has_T_405 ? 64'hffffffffffffffff : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [63:0] _rmask_T_140 = _has_T_407 ? 64'hffffffffffffffff : _rmask_T_138; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [63:0] _rmask_T_142 = _has_T_409 ? 64'hffffffffffffffff : _rmask_T_140; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [63:0] _rmask_T_144 = _has_T_411 ? 64'hffffffffffffffff : _rmask_T_142; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [63:0] _rmask_T_146 = _has_T_413 ? 64'hffffffffffffffff : _rmask_T_144; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [63:0] _rmask_T_148 = _has_T_415 ? 64'hffffffffffffffff : _rmask_T_146; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [63:0] _rmask_T_150 = _has_T_417 ? 64'hffffffffffffffff : _rmask_T_148; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [63:0] _rmask_T_152 = _has_T_419 ? 64'hffffffffffffffff : _rmask_T_150; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [63:0] _rmask_T_154 = _has_T_421 ? 64'hffffffffffffffff : _rmask_T_152; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [63:0] _rmask_T_156 = _has_T_423 ? 64'hffffffffffffffff : _rmask_T_154; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [63:0] _rmask_T_158 = _has_T_425 ? 64'hffffffffffffffff : _rmask_T_156; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [63:0] _rmask_T_160 = _has_T_427 ? 64'hffffffffffffffff : _rmask_T_158; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [63:0] _rmask_T_162 = _has_T_429 ? 64'hffffffffffffffff : _rmask_T_160; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [63:0] rmask_3 = _has_T_431 ? 64'hffffffffffffffff : _rmask_T_162; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 25:44]
  wire [63:0] _GEN_11246 = {{32'd0}, nowCSR_3[31:0]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 32:40]
  wire [63:0] _rData_T_37 = _GEN_11246 & rmask_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 32:40]
  wire [63:0] _GEN_10800 = has_15 ? _rData_T_37 : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 31:17 32:15 35:15]
  wire [63:0] _GEN_10801 = io_now_csr_IALIGN == 8'h20 ? {{32'd0}, _rData_T_41} : _GEN_10800; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:46 46:19]
  wire [63:0] _GEN_10802 = _has_T_427 ? _GEN_10801 : _GEN_10800; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire [63:0] _rData_T_47 = 64'hfffffffffffffffc & io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 46:63]
  wire [63:0] _rData_T_43 = nowCSR_3 & rmask_3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 32:40]
  wire [63:0] _GEN_10803 = has_15 ? _rData_T_43 : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 31:17 32:15 35:15]
  wire [63:0] _GEN_10804 = io_now_csr_IALIGN == 8'h20 ? _rData_T_47 : _GEN_10803; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 45:46 46:19]
  wire [63:0] _GEN_10805 = _has_T_427 ? _GEN_10804 : _GEN_10803; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 39:20]
  wire [63:0] _GEN_10806 = _T_1846 ? _GEN_10805 : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 27:25 52:27]
  wire [63:0] rData_3 = _T_1829 ? _GEN_10802 : _GEN_10806; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 52:27]
  wire [63:0] _T_1802 = {59'h0,rs1}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [63:0] _T_1803 = ~_T_1802; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:63]
  wire [63:0] _T_1804 = rData_3 & _T_1803; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 142:61]
  wire [63:0] _T_1761 = rData_3 | _T_1802; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 131:61]
  wire [63:0] _T_1683 = ~_GEN_101; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:63]
  wire [63:0] _T_1684 = rData_3 & _T_1683; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 110:61]
  wire [63:0] _T_1642 = rData_3 | _GEN_101; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 99:61]
  wire [63:0] _GEN_9915 = csrAddr == 12'h341 ? _GEN_101 : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_9925 = has_15 ? _GEN_9915 : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [63:0] _GEN_9969 = _T_1793 ? _GEN_9925 : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_10023 = _T_1592 ? _GEN_9969 : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10083 = csrAddr == 12'h341 ? _T_1642 : _GEN_10023; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10093 = has_15 ? _GEN_10083 : _GEN_10023; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10105 = _T_1794 ? _GEN_10093 : _GEN_10023; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [63:0] _GEN_10149 = _T_1751 ? _GEN_10105 : _GEN_10023; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10203 = _T_1625 ? _GEN_10149 : _GEN_10023; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10263 = csrAddr == 12'h341 ? _T_1684 : _GEN_10203; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10273 = has_15 ? _GEN_10263 : _GEN_10203; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10285 = _T_1794 ? _GEN_10273 : _GEN_10203; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [63:0] _GEN_10329 = _T_1793 ? _GEN_10285 : _GEN_10203; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10383 = _T_1667 ? _GEN_10329 : _GEN_10203; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10467 = csrAddr == 12'h341 ? _T_1802 : _GEN_10383; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10477 = has_15 ? _GEN_10467 : _GEN_10383; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10521 = _T_1793 ? _GEN_10477 : _GEN_10383; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10575 = _T_1709 ? _GEN_10521 : _GEN_10383; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10635 = csrAddr == 12'h341 ? _T_1761 : _GEN_10575; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10645 = has_15 ? _GEN_10635 : _GEN_10575; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10657 = _T_1794 ? _GEN_10645 : _GEN_10575; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [63:0] _GEN_10701 = ~isIllegalWrite_4 ? _GEN_10657 : _GEN_10575; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10755 = _T_1743 ? _GEN_10701 : _GEN_10575; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10815 = csrAddr == 12'h341 ? _T_1804 : _GEN_10755; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10825 = has_15 ? _GEN_10815 : _GEN_10755; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10837 = rs1 != 5'h0 ? _GEN_10825 : _GEN_10755; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [63:0] _GEN_10881 = ~isIllegalWrite_5 ? _GEN_10837 : _GEN_10755; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10935 = _T_1786 ? _GEN_10881 : _GEN_10755; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_11008 = _T_1846 ? io_now_pc : _GEN_10935; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 186:35]
  wire [63:0] _GEN_11018 = _T_1829 ? io_now_pc : _GEN_11008; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 186:35]
  wire [63:0] _GEN_11042 = delegS ? _GEN_10935 : _GEN_11018; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [63:0] _GEN_11056 = raiseExceptionIntr ? _GEN_11042 : _GEN_10935; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [1:0] _GEN_9799 = io_now_internal_privilegeMode == 2'h3 ? next_reg_mstatusStruct_10_mpp : _GEN_9794; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 88:48 92:35]
  wire [63:0] _GEN_9800 = io_now_internal_privilegeMode == 2'h3 ? _next_csr_mstatus_T_1 : _GEN_9795; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 100:24 88:48]
  wire  _GEN_9802 = io_now_internal_privilegeMode == 2'h3 | _GEN_9797; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 103:25 88:48]
  wire [63:0] _GEN_9803 = io_now_internal_privilegeMode == 2'h3 ? io_now_csr_mepc : _GEN_9798; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 104:25 88:48]
  wire [1:0] _GEN_9813 = _T_1573 ? _GEN_9799 : _GEN_9794; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [63:0] _GEN_9814 = _T_1573 ? _GEN_9800 : _GEN_9795; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire  _GEN_9816 = _T_1573 ? _GEN_9802 : _GEN_9797; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire [63:0] _GEN_9817 = _T_1573 ? _GEN_9803 : _GEN_9798; // @[src/main/scala/rvspeccore/core/spec/instset/Privileged.scala 56:22]
  wire  _T_1600 = rd != 5'h0; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:17]
  wire [63:0] _GEN_9845 = 5'h1 == rd ? rData_3 : _GEN_9743; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9846 = 5'h2 == rd ? rData_3 : _GEN_9744; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9847 = 5'h3 == rd ? rData_3 : _GEN_9745; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9848 = 5'h4 == rd ? rData_3 : _GEN_9746; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9849 = 5'h5 == rd ? rData_3 : _GEN_9747; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9850 = 5'h6 == rd ? rData_3 : _GEN_9748; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9851 = 5'h7 == rd ? rData_3 : _GEN_9749; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9852 = 5'h8 == rd ? rData_3 : _GEN_9750; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9853 = 5'h9 == rd ? rData_3 : _GEN_9751; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9854 = 5'ha == rd ? rData_3 : _GEN_9752; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9855 = 5'hb == rd ? rData_3 : _GEN_9753; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9856 = 5'hc == rd ? rData_3 : _GEN_9754; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9857 = 5'hd == rd ? rData_3 : _GEN_9755; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9858 = 5'he == rd ? rData_3 : _GEN_9756; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9859 = 5'hf == rd ? rData_3 : _GEN_9757; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9860 = 5'h10 == rd ? rData_3 : _GEN_9758; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9861 = 5'h11 == rd ? rData_3 : _GEN_9759; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9862 = 5'h12 == rd ? rData_3 : _GEN_9760; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9863 = 5'h13 == rd ? rData_3 : _GEN_9761; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9864 = 5'h14 == rd ? rData_3 : _GEN_9762; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9865 = 5'h15 == rd ? rData_3 : _GEN_9763; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9866 = 5'h16 == rd ? rData_3 : _GEN_9764; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9867 = 5'h17 == rd ? rData_3 : _GEN_9765; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9868 = 5'h18 == rd ? rData_3 : _GEN_9766; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9869 = 5'h19 == rd ? rData_3 : _GEN_9767; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9870 = 5'h1a == rd ? rData_3 : _GEN_9768; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9871 = 5'h1b == rd ? rData_3 : _GEN_9769; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9872 = 5'h1c == rd ? rData_3 : _GEN_9770; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9873 = 5'h1d == rd ? rData_3 : _GEN_9771; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9874 = 5'h1e == rd ? rData_3 : _GEN_9772; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9875 = 5'h1f == rd ? rData_3 : _GEN_9773; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 87:{24,24}]
  wire [63:0] _GEN_9877 = rd != 5'h0 ? _GEN_9845 : _GEN_9743; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9878 = rd != 5'h0 ? _GEN_9846 : _GEN_9744; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9879 = rd != 5'h0 ? _GEN_9847 : _GEN_9745; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9880 = rd != 5'h0 ? _GEN_9848 : _GEN_9746; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9881 = rd != 5'h0 ? _GEN_9849 : _GEN_9747; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9882 = rd != 5'h0 ? _GEN_9850 : _GEN_9748; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9883 = rd != 5'h0 ? _GEN_9851 : _GEN_9749; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9884 = rd != 5'h0 ? _GEN_9852 : _GEN_9750; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9885 = rd != 5'h0 ? _GEN_9853 : _GEN_9751; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9886 = rd != 5'h0 ? _GEN_9854 : _GEN_9752; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9887 = rd != 5'h0 ? _GEN_9855 : _GEN_9753; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9888 = rd != 5'h0 ? _GEN_9856 : _GEN_9754; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9889 = rd != 5'h0 ? _GEN_9857 : _GEN_9755; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9890 = rd != 5'h0 ? _GEN_9858 : _GEN_9756; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9891 = rd != 5'h0 ? _GEN_9859 : _GEN_9757; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9892 = rd != 5'h0 ? _GEN_9860 : _GEN_9758; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9893 = rd != 5'h0 ? _GEN_9861 : _GEN_9759; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9894 = rd != 5'h0 ? _GEN_9862 : _GEN_9760; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9895 = rd != 5'h0 ? _GEN_9863 : _GEN_9761; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9896 = rd != 5'h0 ? _GEN_9864 : _GEN_9762; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9897 = rd != 5'h0 ? _GEN_9865 : _GEN_9763; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9898 = rd != 5'h0 ? _GEN_9866 : _GEN_9764; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9899 = rd != 5'h0 ? _GEN_9867 : _GEN_9765; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9900 = rd != 5'h0 ? _GEN_9868 : _GEN_9766; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9901 = rd != 5'h0 ? _GEN_9869 : _GEN_9767; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9902 = rd != 5'h0 ? _GEN_9870 : _GEN_9768; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9903 = rd != 5'h0 ? _GEN_9871 : _GEN_9769; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9904 = rd != 5'h0 ? _GEN_9872 : _GEN_9770; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9905 = rd != 5'h0 ? _GEN_9873 : _GEN_9771; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9906 = rd != 5'h0 ? _GEN_9874 : _GEN_9772; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9907 = rd != 5'h0 ? _GEN_9875 : _GEN_9773; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 86:26]
  wire [63:0] _GEN_9908 = csrAddr == 12'h301 ? _GEN_101 : io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  next_csr_mstatus_mstatusOld_pad4 = _GEN_101[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_sie = _GEN_101[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_pad3 = _GEN_101[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_mie = _GEN_101[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_pad2 = _GEN_101[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_spie = _GEN_101[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_ube = _GEN_101[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_mpie = _GEN_101[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_spp = _GEN_101[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_vs = _GEN_101[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_mpp = _GEN_101[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_fs = _GEN_101[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_xs = _GEN_101[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_mprv = _GEN_101[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_sum = _GEN_101[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_mxr = _GEN_101[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_tvm = _GEN_101[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_tw = _GEN_101[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_tsr = _GEN_101[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [8:0] next_csr_mstatus_mstatusOld_pad0 = _GEN_101[31:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_uxl = _GEN_101[33:32]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_sxl = _GEN_101[35:34]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_sbe = _GEN_101[36]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_mbe = _GEN_101[37]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [24:0] next_csr_mstatus_mstatusOld_pad1 = _GEN_101[62:38]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_sd = _GEN_101[63]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [5:0] next_csr_mstatus_mstatusNew_lo_lo = {next_csr_mstatus_mstatusOld_spie,next_csr_mstatus_mstatusOld_pad2,
    next_csr_mstatus_mstatusOld_mie,next_csr_mstatus_mstatusOld_pad3,next_csr_mstatus_mstatusOld_sie,
    next_csr_mstatus_mstatusOld_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [16:0] next_csr_mstatus_mstatusNew_lo = {next_csr_mstatus_mstatusOld_xs,next_csr_mstatus_mstatusOld_fs,
    next_csr_mstatus_mstatusOld_mpp,next_csr_mstatus_mstatusOld_vs,next_csr_mstatus_mstatusOld_spp,
    next_csr_mstatus_mstatusOld_mpie,next_csr_mstatus_mstatusOld_ube,next_csr_mstatus_mstatusNew_lo_lo}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [5:0] next_csr_mstatus_mstatusNew_hi_lo = {next_csr_mstatus_mstatusOld_tsr,next_csr_mstatus_mstatusOld_tw,
    next_csr_mstatus_mstatusOld_tvm,next_csr_mstatus_mstatusOld_mxr,next_csr_mstatus_mstatusOld_sum,
    next_csr_mstatus_mstatusOld_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [63:0] _next_csr_mstatus_mstatusNew_T_1 = {next_csr_mstatus_mstatusOld_sd,next_csr_mstatus_mstatusOld_pad1,
    next_csr_mstatus_mstatusOld_mbe,next_csr_mstatus_mstatusOld_sbe,next_csr_mstatus_mstatusOld_sxl,
    next_csr_mstatus_mstatusOld_uxl,next_csr_mstatus_mstatusOld_pad0,next_csr_mstatus_mstatusNew_hi_lo,
    next_csr_mstatus_mstatusNew_lo}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [63:0] next_csr_mstatus_mstatusNew = {next_csr_mstatus_mstatusOld_fs == 2'h3,_next_csr_mstatus_mstatusNew_T_1[62:
    0]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:27]
  wire [63:0] _GEN_9909 = csrAddr == 12'h300 ? next_csr_mstatus_mstatusNew : _GEN_9814; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_9910 = csrAddr == 12'h340 ? _GEN_101 : io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_9911 = csrAddr == 12'h305 ? _GEN_101 : io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_9912 = csrAddr == 12'h306 ? _GEN_101 : io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _next_csr_mip_T_1 = io_now_csr_mip & 64'h80; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:51]
  wire [63:0] _next_csr_mip_T_2 = _GEN_101 & 64'h77f; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:80]
  wire [63:0] _next_csr_mip_T_3 = _next_csr_mip_T_1 | _next_csr_mip_T_2; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:72]
  wire [63:0] _GEN_9913 = csrAddr == 12'h344 ? _next_csr_mip_T_3 : io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_9914 = csrAddr == 12'h304 ? _GEN_101 : io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_9916 = csrAddr == 12'h342 ? _GEN_101 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_9917 = csrAddr == 12'h343 ? _GEN_101 : _GEN_1995; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_9918 = has_15 ? _GEN_9908 : io_now_csr_misa; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [63:0] _GEN_9919 = has_15 ? _GEN_9909 : _GEN_9814; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_9920 = has_15 ? _GEN_9910 : io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [63:0] _GEN_9921 = has_15 ? _GEN_9911 : io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [63:0] _GEN_9922 = has_15 ? _GEN_9912 : io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [63:0] _GEN_9923 = has_15 ? _GEN_9913 : io_now_csr_mip; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [63:0] _GEN_9924 = has_15 ? _GEN_9914 : io_now_csr_mie; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [63:0] _GEN_9926 = has_15 ? _GEN_9916 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [63:0] _GEN_9927 = has_15 ? _GEN_9917 : _GEN_1995; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_9931 = _T_1793 ? _GEN_9877 : _GEN_9743; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9932 = _T_1793 ? _GEN_9878 : _GEN_9744; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9933 = _T_1793 ? _GEN_9879 : _GEN_9745; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9934 = _T_1793 ? _GEN_9880 : _GEN_9746; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9935 = _T_1793 ? _GEN_9881 : _GEN_9747; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9936 = _T_1793 ? _GEN_9882 : _GEN_9748; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9937 = _T_1793 ? _GEN_9883 : _GEN_9749; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9938 = _T_1793 ? _GEN_9884 : _GEN_9750; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9939 = _T_1793 ? _GEN_9885 : _GEN_9751; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9940 = _T_1793 ? _GEN_9886 : _GEN_9752; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9941 = _T_1793 ? _GEN_9887 : _GEN_9753; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9942 = _T_1793 ? _GEN_9888 : _GEN_9754; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9943 = _T_1793 ? _GEN_9889 : _GEN_9755; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9944 = _T_1793 ? _GEN_9890 : _GEN_9756; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9945 = _T_1793 ? _GEN_9891 : _GEN_9757; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9946 = _T_1793 ? _GEN_9892 : _GEN_9758; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9947 = _T_1793 ? _GEN_9893 : _GEN_9759; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9948 = _T_1793 ? _GEN_9894 : _GEN_9760; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9949 = _T_1793 ? _GEN_9895 : _GEN_9761; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9950 = _T_1793 ? _GEN_9896 : _GEN_9762; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9951 = _T_1793 ? _GEN_9897 : _GEN_9763; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9952 = _T_1793 ? _GEN_9898 : _GEN_9764; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9953 = _T_1793 ? _GEN_9899 : _GEN_9765; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9954 = _T_1793 ? _GEN_9900 : _GEN_9766; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9955 = _T_1793 ? _GEN_9901 : _GEN_9767; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9956 = _T_1793 ? _GEN_9902 : _GEN_9768; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9957 = _T_1793 ? _GEN_9903 : _GEN_9769; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9958 = _T_1793 ? _GEN_9904 : _GEN_9770; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9959 = _T_1793 ? _GEN_9905 : _GEN_9771; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9960 = _T_1793 ? _GEN_9906 : _GEN_9772; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9961 = _T_1793 ? _GEN_9907 : _GEN_9773; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9962 = _T_1793 ? _GEN_9918 : io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9963 = _T_1793 ? _GEN_9919 : _GEN_9814; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9964 = _T_1793 ? _GEN_9920 : io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9965 = _T_1793 ? _GEN_9921 : io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9966 = _T_1793 ? _GEN_9922 : io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9967 = _T_1793 ? _GEN_9923 : io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9968 = _T_1793 ? _GEN_9924 : io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9970 = _T_1793 ? _GEN_9926 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9971 = _T_1793 ? _GEN_9927 : _GEN_1995; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 85:27]
  wire [63:0] _GEN_9985 = _T_1592 ? _GEN_9931 : _GEN_9743; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_9986 = _T_1592 ? _GEN_9932 : _GEN_9744; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_9987 = _T_1592 ? _GEN_9933 : _GEN_9745; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_9988 = _T_1592 ? _GEN_9934 : _GEN_9746; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_9989 = _T_1592 ? _GEN_9935 : _GEN_9747; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_9990 = _T_1592 ? _GEN_9936 : _GEN_9748; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_9991 = _T_1592 ? _GEN_9937 : _GEN_9749; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_9992 = _T_1592 ? _GEN_9938 : _GEN_9750; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_9993 = _T_1592 ? _GEN_9939 : _GEN_9751; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_9994 = _T_1592 ? _GEN_9940 : _GEN_9752; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_9995 = _T_1592 ? _GEN_9941 : _GEN_9753; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_9996 = _T_1592 ? _GEN_9942 : _GEN_9754; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_9997 = _T_1592 ? _GEN_9943 : _GEN_9755; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_9998 = _T_1592 ? _GEN_9944 : _GEN_9756; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_9999 = _T_1592 ? _GEN_9945 : _GEN_9757; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10000 = _T_1592 ? _GEN_9946 : _GEN_9758; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10001 = _T_1592 ? _GEN_9947 : _GEN_9759; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10002 = _T_1592 ? _GEN_9948 : _GEN_9760; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10003 = _T_1592 ? _GEN_9949 : _GEN_9761; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10004 = _T_1592 ? _GEN_9950 : _GEN_9762; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10005 = _T_1592 ? _GEN_9951 : _GEN_9763; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10006 = _T_1592 ? _GEN_9952 : _GEN_9764; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10007 = _T_1592 ? _GEN_9953 : _GEN_9765; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10008 = _T_1592 ? _GEN_9954 : _GEN_9766; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10009 = _T_1592 ? _GEN_9955 : _GEN_9767; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10010 = _T_1592 ? _GEN_9956 : _GEN_9768; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10011 = _T_1592 ? _GEN_9957 : _GEN_9769; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10012 = _T_1592 ? _GEN_9958 : _GEN_9770; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10013 = _T_1592 ? _GEN_9959 : _GEN_9771; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10014 = _T_1592 ? _GEN_9960 : _GEN_9772; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10015 = _T_1592 ? _GEN_9961 : _GEN_9773; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10016 = _T_1592 ? _GEN_9962 : io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10017 = _T_1592 ? _GEN_9963 : _GEN_9814; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10018 = _T_1592 ? _GEN_9964 : io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10019 = _T_1592 ? _GEN_9965 : io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10020 = _T_1592 ? _GEN_9966 : io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10021 = _T_1592 ? _GEN_9967 : io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10022 = _T_1592 ? _GEN_9968 : io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10024 = _T_1592 ? _GEN_9970 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10025 = _T_1592 ? _GEN_9971 : _GEN_1995; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 82:23]
  wire [63:0] _GEN_10037 = 5'h1 == rd ? rData_3 : _GEN_9985; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10038 = 5'h2 == rd ? rData_3 : _GEN_9986; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10039 = 5'h3 == rd ? rData_3 : _GEN_9987; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10040 = 5'h4 == rd ? rData_3 : _GEN_9988; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10041 = 5'h5 == rd ? rData_3 : _GEN_9989; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10042 = 5'h6 == rd ? rData_3 : _GEN_9990; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10043 = 5'h7 == rd ? rData_3 : _GEN_9991; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10044 = 5'h8 == rd ? rData_3 : _GEN_9992; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10045 = 5'h9 == rd ? rData_3 : _GEN_9993; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10046 = 5'ha == rd ? rData_3 : _GEN_9994; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10047 = 5'hb == rd ? rData_3 : _GEN_9995; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10048 = 5'hc == rd ? rData_3 : _GEN_9996; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10049 = 5'hd == rd ? rData_3 : _GEN_9997; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10050 = 5'he == rd ? rData_3 : _GEN_9998; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10051 = 5'hf == rd ? rData_3 : _GEN_9999; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10052 = 5'h10 == rd ? rData_3 : _GEN_10000; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10053 = 5'h11 == rd ? rData_3 : _GEN_10001; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10054 = 5'h12 == rd ? rData_3 : _GEN_10002; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10055 = 5'h13 == rd ? rData_3 : _GEN_10003; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10056 = 5'h14 == rd ? rData_3 : _GEN_10004; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10057 = 5'h15 == rd ? rData_3 : _GEN_10005; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10058 = 5'h16 == rd ? rData_3 : _GEN_10006; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10059 = 5'h17 == rd ? rData_3 : _GEN_10007; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10060 = 5'h18 == rd ? rData_3 : _GEN_10008; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10061 = 5'h19 == rd ? rData_3 : _GEN_10009; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10062 = 5'h1a == rd ? rData_3 : _GEN_10010; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10063 = 5'h1b == rd ? rData_3 : _GEN_10011; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10064 = 5'h1c == rd ? rData_3 : _GEN_10012; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10065 = 5'h1d == rd ? rData_3 : _GEN_10013; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10066 = 5'h1e == rd ? rData_3 : _GEN_10014; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10067 = 5'h1f == rd ? rData_3 : _GEN_10015; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 97:{22,22}]
  wire [63:0] _GEN_10076 = csrAddr == 12'h301 ? _T_1642 : _GEN_10016; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  next_csr_mstatus_mstatusOld_1_pad4 = _T_1642[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_sie = _T_1642[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_pad3 = _T_1642[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_mie = _T_1642[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_pad2 = _T_1642[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_spie = _T_1642[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_ube = _T_1642[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_mpie = _T_1642[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_spp = _T_1642[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_1_vs = _T_1642[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_1_mpp = _T_1642[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_1_fs = _T_1642[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_1_xs = _T_1642[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_mprv = _T_1642[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_sum = _T_1642[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_mxr = _T_1642[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_tvm = _T_1642[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_tw = _T_1642[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_tsr = _T_1642[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [8:0] next_csr_mstatus_mstatusOld_1_pad0 = _T_1642[31:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_1_uxl = _T_1642[33:32]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_1_sxl = _T_1642[35:34]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_sbe = _T_1642[36]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_mbe = _T_1642[37]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [24:0] next_csr_mstatus_mstatusOld_1_pad1 = _T_1642[62:38]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_1_sd = _T_1642[63]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [5:0] next_csr_mstatus_mstatusNew_lo_lo_1 = {next_csr_mstatus_mstatusOld_1_spie,
    next_csr_mstatus_mstatusOld_1_pad2,next_csr_mstatus_mstatusOld_1_mie,next_csr_mstatus_mstatusOld_1_pad3,
    next_csr_mstatus_mstatusOld_1_sie,next_csr_mstatus_mstatusOld_1_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [16:0] next_csr_mstatus_mstatusNew_lo_1 = {next_csr_mstatus_mstatusOld_1_xs,next_csr_mstatus_mstatusOld_1_fs,
    next_csr_mstatus_mstatusOld_1_mpp,next_csr_mstatus_mstatusOld_1_vs,next_csr_mstatus_mstatusOld_1_spp,
    next_csr_mstatus_mstatusOld_1_mpie,next_csr_mstatus_mstatusOld_1_ube,next_csr_mstatus_mstatusNew_lo_lo_1}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [5:0] next_csr_mstatus_mstatusNew_hi_lo_1 = {next_csr_mstatus_mstatusOld_1_tsr,next_csr_mstatus_mstatusOld_1_tw,
    next_csr_mstatus_mstatusOld_1_tvm,next_csr_mstatus_mstatusOld_1_mxr,next_csr_mstatus_mstatusOld_1_sum,
    next_csr_mstatus_mstatusOld_1_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [63:0] _next_csr_mstatus_mstatusNew_T_4 = {next_csr_mstatus_mstatusOld_1_sd,next_csr_mstatus_mstatusOld_1_pad1,
    next_csr_mstatus_mstatusOld_1_mbe,next_csr_mstatus_mstatusOld_1_sbe,next_csr_mstatus_mstatusOld_1_sxl,
    next_csr_mstatus_mstatusOld_1_uxl,next_csr_mstatus_mstatusOld_1_pad0,next_csr_mstatus_mstatusNew_hi_lo_1,
    next_csr_mstatus_mstatusNew_lo_1}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [63:0] next_csr_mstatus_mstatusNew_1 = {next_csr_mstatus_mstatusOld_1_fs == 2'h3,_next_csr_mstatus_mstatusNew_T_4
    [62:0]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:27]
  wire [63:0] _GEN_10077 = csrAddr == 12'h300 ? next_csr_mstatus_mstatusNew_1 : _GEN_10017; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10078 = csrAddr == 12'h340 ? _T_1642 : _GEN_10018; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10079 = csrAddr == 12'h305 ? _T_1642 : _GEN_10019; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10080 = csrAddr == 12'h306 ? _T_1642 : _GEN_10020; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _next_csr_mip_T_6 = _T_1642 & 64'h77f; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:80]
  wire [63:0] _next_csr_mip_T_7 = _next_csr_mip_T_1 | _next_csr_mip_T_6; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:72]
  wire [63:0] _GEN_10081 = csrAddr == 12'h344 ? _next_csr_mip_T_7 : _GEN_10021; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10082 = csrAddr == 12'h304 ? _T_1642 : _GEN_10022; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10084 = csrAddr == 12'h342 ? _T_1642 : _GEN_10024; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10085 = csrAddr == 12'h343 ? _T_1642 : _GEN_10025; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10086 = has_15 ? _GEN_10076 : _GEN_10016; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10087 = has_15 ? _GEN_10077 : _GEN_10017; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10088 = has_15 ? _GEN_10078 : _GEN_10018; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10089 = has_15 ? _GEN_10079 : _GEN_10019; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10090 = has_15 ? _GEN_10080 : _GEN_10020; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10091 = has_15 ? _GEN_10081 : _GEN_10021; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10092 = has_15 ? _GEN_10082 : _GEN_10022; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10094 = has_15 ? _GEN_10084 : _GEN_10024; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10095 = has_15 ? _GEN_10085 : _GEN_10025; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10098 = _T_1794 ? _GEN_10086 : _GEN_10016; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [63:0] _GEN_10099 = _T_1794 ? _GEN_10087 : _GEN_10017; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [63:0] _GEN_10100 = _T_1794 ? _GEN_10088 : _GEN_10018; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [63:0] _GEN_10101 = _T_1794 ? _GEN_10089 : _GEN_10019; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [63:0] _GEN_10102 = _T_1794 ? _GEN_10090 : _GEN_10020; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [63:0] _GEN_10103 = _T_1794 ? _GEN_10091 : _GEN_10021; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [63:0] _GEN_10104 = _T_1794 ? _GEN_10092 : _GEN_10022; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [63:0] _GEN_10106 = _T_1794 ? _GEN_10094 : _GEN_10024; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [63:0] _GEN_10107 = _T_1794 ? _GEN_10095 : _GEN_10025; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 98:27]
  wire [63:0] _GEN_10111 = _T_1751 ? _GEN_10037 : _GEN_9985; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10112 = _T_1751 ? _GEN_10038 : _GEN_9986; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10113 = _T_1751 ? _GEN_10039 : _GEN_9987; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10114 = _T_1751 ? _GEN_10040 : _GEN_9988; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10115 = _T_1751 ? _GEN_10041 : _GEN_9989; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10116 = _T_1751 ? _GEN_10042 : _GEN_9990; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10117 = _T_1751 ? _GEN_10043 : _GEN_9991; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10118 = _T_1751 ? _GEN_10044 : _GEN_9992; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10119 = _T_1751 ? _GEN_10045 : _GEN_9993; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10120 = _T_1751 ? _GEN_10046 : _GEN_9994; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10121 = _T_1751 ? _GEN_10047 : _GEN_9995; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10122 = _T_1751 ? _GEN_10048 : _GEN_9996; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10123 = _T_1751 ? _GEN_10049 : _GEN_9997; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10124 = _T_1751 ? _GEN_10050 : _GEN_9998; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10125 = _T_1751 ? _GEN_10051 : _GEN_9999; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10126 = _T_1751 ? _GEN_10052 : _GEN_10000; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10127 = _T_1751 ? _GEN_10053 : _GEN_10001; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10128 = _T_1751 ? _GEN_10054 : _GEN_10002; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10129 = _T_1751 ? _GEN_10055 : _GEN_10003; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10130 = _T_1751 ? _GEN_10056 : _GEN_10004; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10131 = _T_1751 ? _GEN_10057 : _GEN_10005; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10132 = _T_1751 ? _GEN_10058 : _GEN_10006; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10133 = _T_1751 ? _GEN_10059 : _GEN_10007; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10134 = _T_1751 ? _GEN_10060 : _GEN_10008; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10135 = _T_1751 ? _GEN_10061 : _GEN_10009; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10136 = _T_1751 ? _GEN_10062 : _GEN_10010; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10137 = _T_1751 ? _GEN_10063 : _GEN_10011; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10138 = _T_1751 ? _GEN_10064 : _GEN_10012; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10139 = _T_1751 ? _GEN_10065 : _GEN_10013; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10140 = _T_1751 ? _GEN_10066 : _GEN_10014; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10141 = _T_1751 ? _GEN_10067 : _GEN_10015; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10142 = _T_1751 ? _GEN_10098 : _GEN_10016; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10143 = _T_1751 ? _GEN_10099 : _GEN_10017; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10144 = _T_1751 ? _GEN_10100 : _GEN_10018; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10145 = _T_1751 ? _GEN_10101 : _GEN_10019; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10146 = _T_1751 ? _GEN_10102 : _GEN_10020; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10147 = _T_1751 ? _GEN_10103 : _GEN_10021; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10148 = _T_1751 ? _GEN_10104 : _GEN_10022; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10150 = _T_1751 ? _GEN_10106 : _GEN_10024; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10151 = _T_1751 ? _GEN_10107 : _GEN_10025; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 96:49]
  wire [63:0] _GEN_10165 = _T_1625 ? _GEN_10111 : _GEN_9985; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10166 = _T_1625 ? _GEN_10112 : _GEN_9986; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10167 = _T_1625 ? _GEN_10113 : _GEN_9987; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10168 = _T_1625 ? _GEN_10114 : _GEN_9988; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10169 = _T_1625 ? _GEN_10115 : _GEN_9989; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10170 = _T_1625 ? _GEN_10116 : _GEN_9990; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10171 = _T_1625 ? _GEN_10117 : _GEN_9991; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10172 = _T_1625 ? _GEN_10118 : _GEN_9992; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10173 = _T_1625 ? _GEN_10119 : _GEN_9993; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10174 = _T_1625 ? _GEN_10120 : _GEN_9994; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10175 = _T_1625 ? _GEN_10121 : _GEN_9995; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10176 = _T_1625 ? _GEN_10122 : _GEN_9996; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10177 = _T_1625 ? _GEN_10123 : _GEN_9997; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10178 = _T_1625 ? _GEN_10124 : _GEN_9998; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10179 = _T_1625 ? _GEN_10125 : _GEN_9999; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10180 = _T_1625 ? _GEN_10126 : _GEN_10000; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10181 = _T_1625 ? _GEN_10127 : _GEN_10001; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10182 = _T_1625 ? _GEN_10128 : _GEN_10002; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10183 = _T_1625 ? _GEN_10129 : _GEN_10003; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10184 = _T_1625 ? _GEN_10130 : _GEN_10004; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10185 = _T_1625 ? _GEN_10131 : _GEN_10005; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10186 = _T_1625 ? _GEN_10132 : _GEN_10006; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10187 = _T_1625 ? _GEN_10133 : _GEN_10007; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10188 = _T_1625 ? _GEN_10134 : _GEN_10008; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10189 = _T_1625 ? _GEN_10135 : _GEN_10009; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10190 = _T_1625 ? _GEN_10136 : _GEN_10010; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10191 = _T_1625 ? _GEN_10137 : _GEN_10011; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10192 = _T_1625 ? _GEN_10138 : _GEN_10012; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10193 = _T_1625 ? _GEN_10139 : _GEN_10013; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10194 = _T_1625 ? _GEN_10140 : _GEN_10014; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10195 = _T_1625 ? _GEN_10141 : _GEN_10015; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10196 = _T_1625 ? _GEN_10142 : _GEN_10016; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10197 = _T_1625 ? _GEN_10143 : _GEN_10017; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10198 = _T_1625 ? _GEN_10144 : _GEN_10018; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10199 = _T_1625 ? _GEN_10145 : _GEN_10019; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10200 = _T_1625 ? _GEN_10146 : _GEN_10020; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10201 = _T_1625 ? _GEN_10147 : _GEN_10021; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10202 = _T_1625 ? _GEN_10148 : _GEN_10022; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10204 = _T_1625 ? _GEN_10150 : _GEN_10024; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10205 = _T_1625 ? _GEN_10151 : _GEN_10025; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 93:23]
  wire [63:0] _GEN_10217 = 5'h1 == rd ? rData_3 : _GEN_10165; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10218 = 5'h2 == rd ? rData_3 : _GEN_10166; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10219 = 5'h3 == rd ? rData_3 : _GEN_10167; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10220 = 5'h4 == rd ? rData_3 : _GEN_10168; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10221 = 5'h5 == rd ? rData_3 : _GEN_10169; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10222 = 5'h6 == rd ? rData_3 : _GEN_10170; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10223 = 5'h7 == rd ? rData_3 : _GEN_10171; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10224 = 5'h8 == rd ? rData_3 : _GEN_10172; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10225 = 5'h9 == rd ? rData_3 : _GEN_10173; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10226 = 5'ha == rd ? rData_3 : _GEN_10174; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10227 = 5'hb == rd ? rData_3 : _GEN_10175; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10228 = 5'hc == rd ? rData_3 : _GEN_10176; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10229 = 5'hd == rd ? rData_3 : _GEN_10177; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10230 = 5'he == rd ? rData_3 : _GEN_10178; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10231 = 5'hf == rd ? rData_3 : _GEN_10179; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10232 = 5'h10 == rd ? rData_3 : _GEN_10180; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10233 = 5'h11 == rd ? rData_3 : _GEN_10181; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10234 = 5'h12 == rd ? rData_3 : _GEN_10182; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10235 = 5'h13 == rd ? rData_3 : _GEN_10183; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10236 = 5'h14 == rd ? rData_3 : _GEN_10184; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10237 = 5'h15 == rd ? rData_3 : _GEN_10185; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10238 = 5'h16 == rd ? rData_3 : _GEN_10186; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10239 = 5'h17 == rd ? rData_3 : _GEN_10187; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10240 = 5'h18 == rd ? rData_3 : _GEN_10188; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10241 = 5'h19 == rd ? rData_3 : _GEN_10189; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10242 = 5'h1a == rd ? rData_3 : _GEN_10190; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10243 = 5'h1b == rd ? rData_3 : _GEN_10191; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10244 = 5'h1c == rd ? rData_3 : _GEN_10192; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10245 = 5'h1d == rd ? rData_3 : _GEN_10193; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10246 = 5'h1e == rd ? rData_3 : _GEN_10194; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10247 = 5'h1f == rd ? rData_3 : _GEN_10195; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 107:{22,22}]
  wire [63:0] _GEN_10256 = csrAddr == 12'h301 ? _T_1684 : _GEN_10196; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  next_csr_mstatus_mstatusOld_2_pad4 = _T_1684[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_sie = _T_1684[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_pad3 = _T_1684[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_mie = _T_1684[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_pad2 = _T_1684[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_spie = _T_1684[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_ube = _T_1684[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_mpie = _T_1684[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_spp = _T_1684[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_2_vs = _T_1684[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_2_mpp = _T_1684[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_2_fs = _T_1684[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_2_xs = _T_1684[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_mprv = _T_1684[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_sum = _T_1684[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_mxr = _T_1684[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_tvm = _T_1684[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_tw = _T_1684[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_tsr = _T_1684[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [8:0] next_csr_mstatus_mstatusOld_2_pad0 = _T_1684[31:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_2_uxl = _T_1684[33:32]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_2_sxl = _T_1684[35:34]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_sbe = _T_1684[36]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_mbe = _T_1684[37]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [24:0] next_csr_mstatus_mstatusOld_2_pad1 = _T_1684[62:38]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_2_sd = _T_1684[63]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [5:0] next_csr_mstatus_mstatusNew_lo_lo_2 = {next_csr_mstatus_mstatusOld_2_spie,
    next_csr_mstatus_mstatusOld_2_pad2,next_csr_mstatus_mstatusOld_2_mie,next_csr_mstatus_mstatusOld_2_pad3,
    next_csr_mstatus_mstatusOld_2_sie,next_csr_mstatus_mstatusOld_2_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [16:0] next_csr_mstatus_mstatusNew_lo_2 = {next_csr_mstatus_mstatusOld_2_xs,next_csr_mstatus_mstatusOld_2_fs,
    next_csr_mstatus_mstatusOld_2_mpp,next_csr_mstatus_mstatusOld_2_vs,next_csr_mstatus_mstatusOld_2_spp,
    next_csr_mstatus_mstatusOld_2_mpie,next_csr_mstatus_mstatusOld_2_ube,next_csr_mstatus_mstatusNew_lo_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [5:0] next_csr_mstatus_mstatusNew_hi_lo_2 = {next_csr_mstatus_mstatusOld_2_tsr,next_csr_mstatus_mstatusOld_2_tw,
    next_csr_mstatus_mstatusOld_2_tvm,next_csr_mstatus_mstatusOld_2_mxr,next_csr_mstatus_mstatusOld_2_sum,
    next_csr_mstatus_mstatusOld_2_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [63:0] _next_csr_mstatus_mstatusNew_T_7 = {next_csr_mstatus_mstatusOld_2_sd,next_csr_mstatus_mstatusOld_2_pad1,
    next_csr_mstatus_mstatusOld_2_mbe,next_csr_mstatus_mstatusOld_2_sbe,next_csr_mstatus_mstatusOld_2_sxl,
    next_csr_mstatus_mstatusOld_2_uxl,next_csr_mstatus_mstatusOld_2_pad0,next_csr_mstatus_mstatusNew_hi_lo_2,
    next_csr_mstatus_mstatusNew_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [63:0] next_csr_mstatus_mstatusNew_2 = {next_csr_mstatus_mstatusOld_2_fs == 2'h3,_next_csr_mstatus_mstatusNew_T_7
    [62:0]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:27]
  wire [63:0] _GEN_10257 = csrAddr == 12'h300 ? next_csr_mstatus_mstatusNew_2 : _GEN_10197; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10258 = csrAddr == 12'h340 ? _T_1684 : _GEN_10198; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10259 = csrAddr == 12'h305 ? _T_1684 : _GEN_10199; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10260 = csrAddr == 12'h306 ? _T_1684 : _GEN_10200; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _next_csr_mip_T_10 = _T_1684 & 64'h77f; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:80]
  wire [63:0] _next_csr_mip_T_11 = _next_csr_mip_T_1 | _next_csr_mip_T_10; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:72]
  wire [63:0] _GEN_10261 = csrAddr == 12'h344 ? _next_csr_mip_T_11 : _GEN_10201; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10262 = csrAddr == 12'h304 ? _T_1684 : _GEN_10202; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10264 = csrAddr == 12'h342 ? _T_1684 : _GEN_10204; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10265 = csrAddr == 12'h343 ? _T_1684 : _GEN_10205; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10266 = has_15 ? _GEN_10256 : _GEN_10196; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10267 = has_15 ? _GEN_10257 : _GEN_10197; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10268 = has_15 ? _GEN_10258 : _GEN_10198; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10269 = has_15 ? _GEN_10259 : _GEN_10199; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10270 = has_15 ? _GEN_10260 : _GEN_10200; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10271 = has_15 ? _GEN_10261 : _GEN_10201; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10272 = has_15 ? _GEN_10262 : _GEN_10202; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10274 = has_15 ? _GEN_10264 : _GEN_10204; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10275 = has_15 ? _GEN_10265 : _GEN_10205; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10278 = _T_1794 ? _GEN_10266 : _GEN_10196; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [63:0] _GEN_10279 = _T_1794 ? _GEN_10267 : _GEN_10197; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [63:0] _GEN_10280 = _T_1794 ? _GEN_10268 : _GEN_10198; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [63:0] _GEN_10281 = _T_1794 ? _GEN_10269 : _GEN_10199; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [63:0] _GEN_10282 = _T_1794 ? _GEN_10270 : _GEN_10200; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [63:0] _GEN_10283 = _T_1794 ? _GEN_10271 : _GEN_10201; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [63:0] _GEN_10284 = _T_1794 ? _GEN_10272 : _GEN_10202; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [63:0] _GEN_10286 = _T_1794 ? _GEN_10274 : _GEN_10204; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [63:0] _GEN_10287 = _T_1794 ? _GEN_10275 : _GEN_10205; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 108:27]
  wire [63:0] _GEN_10291 = _T_1793 ? _GEN_10217 : _GEN_10165; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10292 = _T_1793 ? _GEN_10218 : _GEN_10166; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10293 = _T_1793 ? _GEN_10219 : _GEN_10167; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10294 = _T_1793 ? _GEN_10220 : _GEN_10168; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10295 = _T_1793 ? _GEN_10221 : _GEN_10169; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10296 = _T_1793 ? _GEN_10222 : _GEN_10170; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10297 = _T_1793 ? _GEN_10223 : _GEN_10171; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10298 = _T_1793 ? _GEN_10224 : _GEN_10172; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10299 = _T_1793 ? _GEN_10225 : _GEN_10173; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10300 = _T_1793 ? _GEN_10226 : _GEN_10174; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10301 = _T_1793 ? _GEN_10227 : _GEN_10175; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10302 = _T_1793 ? _GEN_10228 : _GEN_10176; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10303 = _T_1793 ? _GEN_10229 : _GEN_10177; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10304 = _T_1793 ? _GEN_10230 : _GEN_10178; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10305 = _T_1793 ? _GEN_10231 : _GEN_10179; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10306 = _T_1793 ? _GEN_10232 : _GEN_10180; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10307 = _T_1793 ? _GEN_10233 : _GEN_10181; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10308 = _T_1793 ? _GEN_10234 : _GEN_10182; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10309 = _T_1793 ? _GEN_10235 : _GEN_10183; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10310 = _T_1793 ? _GEN_10236 : _GEN_10184; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10311 = _T_1793 ? _GEN_10237 : _GEN_10185; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10312 = _T_1793 ? _GEN_10238 : _GEN_10186; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10313 = _T_1793 ? _GEN_10239 : _GEN_10187; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10314 = _T_1793 ? _GEN_10240 : _GEN_10188; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10315 = _T_1793 ? _GEN_10241 : _GEN_10189; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10316 = _T_1793 ? _GEN_10242 : _GEN_10190; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10317 = _T_1793 ? _GEN_10243 : _GEN_10191; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10318 = _T_1793 ? _GEN_10244 : _GEN_10192; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10319 = _T_1793 ? _GEN_10245 : _GEN_10193; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10320 = _T_1793 ? _GEN_10246 : _GEN_10194; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10321 = _T_1793 ? _GEN_10247 : _GEN_10195; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10322 = _T_1793 ? _GEN_10278 : _GEN_10196; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10323 = _T_1793 ? _GEN_10279 : _GEN_10197; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10324 = _T_1793 ? _GEN_10280 : _GEN_10198; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10325 = _T_1793 ? _GEN_10281 : _GEN_10199; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10326 = _T_1793 ? _GEN_10282 : _GEN_10200; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10327 = _T_1793 ? _GEN_10283 : _GEN_10201; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10328 = _T_1793 ? _GEN_10284 : _GEN_10202; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10330 = _T_1793 ? _GEN_10286 : _GEN_10204; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10331 = _T_1793 ? _GEN_10287 : _GEN_10205; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 106:27]
  wire [63:0] _GEN_10345 = _T_1667 ? _GEN_10291 : _GEN_10165; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10346 = _T_1667 ? _GEN_10292 : _GEN_10166; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10347 = _T_1667 ? _GEN_10293 : _GEN_10167; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10348 = _T_1667 ? _GEN_10294 : _GEN_10168; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10349 = _T_1667 ? _GEN_10295 : _GEN_10169; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10350 = _T_1667 ? _GEN_10296 : _GEN_10170; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10351 = _T_1667 ? _GEN_10297 : _GEN_10171; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10352 = _T_1667 ? _GEN_10298 : _GEN_10172; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10353 = _T_1667 ? _GEN_10299 : _GEN_10173; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10354 = _T_1667 ? _GEN_10300 : _GEN_10174; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10355 = _T_1667 ? _GEN_10301 : _GEN_10175; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10356 = _T_1667 ? _GEN_10302 : _GEN_10176; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10357 = _T_1667 ? _GEN_10303 : _GEN_10177; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10358 = _T_1667 ? _GEN_10304 : _GEN_10178; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10359 = _T_1667 ? _GEN_10305 : _GEN_10179; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10360 = _T_1667 ? _GEN_10306 : _GEN_10180; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10361 = _T_1667 ? _GEN_10307 : _GEN_10181; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10362 = _T_1667 ? _GEN_10308 : _GEN_10182; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10363 = _T_1667 ? _GEN_10309 : _GEN_10183; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10364 = _T_1667 ? _GEN_10310 : _GEN_10184; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10365 = _T_1667 ? _GEN_10311 : _GEN_10185; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10366 = _T_1667 ? _GEN_10312 : _GEN_10186; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10367 = _T_1667 ? _GEN_10313 : _GEN_10187; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10368 = _T_1667 ? _GEN_10314 : _GEN_10188; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10369 = _T_1667 ? _GEN_10315 : _GEN_10189; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10370 = _T_1667 ? _GEN_10316 : _GEN_10190; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10371 = _T_1667 ? _GEN_10317 : _GEN_10191; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10372 = _T_1667 ? _GEN_10318 : _GEN_10192; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10373 = _T_1667 ? _GEN_10319 : _GEN_10193; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10374 = _T_1667 ? _GEN_10320 : _GEN_10194; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10375 = _T_1667 ? _GEN_10321 : _GEN_10195; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10376 = _T_1667 ? _GEN_10322 : _GEN_10196; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10377 = _T_1667 ? _GEN_10323 : _GEN_10197; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10378 = _T_1667 ? _GEN_10324 : _GEN_10198; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10379 = _T_1667 ? _GEN_10325 : _GEN_10199; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10380 = _T_1667 ? _GEN_10326 : _GEN_10200; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10381 = _T_1667 ? _GEN_10327 : _GEN_10201; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10382 = _T_1667 ? _GEN_10328 : _GEN_10202; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10384 = _T_1667 ? _GEN_10330 : _GEN_10204; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10385 = _T_1667 ? _GEN_10331 : _GEN_10205; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 103:23]
  wire [63:0] _GEN_10397 = 5'h1 == rd ? rData_3 : _GEN_10345; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10398 = 5'h2 == rd ? rData_3 : _GEN_10346; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10399 = 5'h3 == rd ? rData_3 : _GEN_10347; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10400 = 5'h4 == rd ? rData_3 : _GEN_10348; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10401 = 5'h5 == rd ? rData_3 : _GEN_10349; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10402 = 5'h6 == rd ? rData_3 : _GEN_10350; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10403 = 5'h7 == rd ? rData_3 : _GEN_10351; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10404 = 5'h8 == rd ? rData_3 : _GEN_10352; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10405 = 5'h9 == rd ? rData_3 : _GEN_10353; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10406 = 5'ha == rd ? rData_3 : _GEN_10354; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10407 = 5'hb == rd ? rData_3 : _GEN_10355; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10408 = 5'hc == rd ? rData_3 : _GEN_10356; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10409 = 5'hd == rd ? rData_3 : _GEN_10357; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10410 = 5'he == rd ? rData_3 : _GEN_10358; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10411 = 5'hf == rd ? rData_3 : _GEN_10359; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10412 = 5'h10 == rd ? rData_3 : _GEN_10360; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10413 = 5'h11 == rd ? rData_3 : _GEN_10361; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10414 = 5'h12 == rd ? rData_3 : _GEN_10362; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10415 = 5'h13 == rd ? rData_3 : _GEN_10363; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10416 = 5'h14 == rd ? rData_3 : _GEN_10364; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10417 = 5'h15 == rd ? rData_3 : _GEN_10365; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10418 = 5'h16 == rd ? rData_3 : _GEN_10366; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10419 = 5'h17 == rd ? rData_3 : _GEN_10367; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10420 = 5'h18 == rd ? rData_3 : _GEN_10368; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10421 = 5'h19 == rd ? rData_3 : _GEN_10369; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10422 = 5'h1a == rd ? rData_3 : _GEN_10370; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10423 = 5'h1b == rd ? rData_3 : _GEN_10371; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10424 = 5'h1c == rd ? rData_3 : _GEN_10372; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10425 = 5'h1d == rd ? rData_3 : _GEN_10373; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10426 = 5'h1e == rd ? rData_3 : _GEN_10374; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10427 = 5'h1f == rd ? rData_3 : _GEN_10375; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 119:{24,24}]
  wire [63:0] _GEN_10429 = _T_1600 ? _GEN_10397 : _GEN_10345; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10430 = _T_1600 ? _GEN_10398 : _GEN_10346; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10431 = _T_1600 ? _GEN_10399 : _GEN_10347; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10432 = _T_1600 ? _GEN_10400 : _GEN_10348; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10433 = _T_1600 ? _GEN_10401 : _GEN_10349; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10434 = _T_1600 ? _GEN_10402 : _GEN_10350; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10435 = _T_1600 ? _GEN_10403 : _GEN_10351; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10436 = _T_1600 ? _GEN_10404 : _GEN_10352; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10437 = _T_1600 ? _GEN_10405 : _GEN_10353; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10438 = _T_1600 ? _GEN_10406 : _GEN_10354; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10439 = _T_1600 ? _GEN_10407 : _GEN_10355; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10440 = _T_1600 ? _GEN_10408 : _GEN_10356; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10441 = _T_1600 ? _GEN_10409 : _GEN_10357; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10442 = _T_1600 ? _GEN_10410 : _GEN_10358; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10443 = _T_1600 ? _GEN_10411 : _GEN_10359; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10444 = _T_1600 ? _GEN_10412 : _GEN_10360; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10445 = _T_1600 ? _GEN_10413 : _GEN_10361; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10446 = _T_1600 ? _GEN_10414 : _GEN_10362; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10447 = _T_1600 ? _GEN_10415 : _GEN_10363; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10448 = _T_1600 ? _GEN_10416 : _GEN_10364; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10449 = _T_1600 ? _GEN_10417 : _GEN_10365; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10450 = _T_1600 ? _GEN_10418 : _GEN_10366; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10451 = _T_1600 ? _GEN_10419 : _GEN_10367; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10452 = _T_1600 ? _GEN_10420 : _GEN_10368; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10453 = _T_1600 ? _GEN_10421 : _GEN_10369; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10454 = _T_1600 ? _GEN_10422 : _GEN_10370; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10455 = _T_1600 ? _GEN_10423 : _GEN_10371; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10456 = _T_1600 ? _GEN_10424 : _GEN_10372; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10457 = _T_1600 ? _GEN_10425 : _GEN_10373; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10458 = _T_1600 ? _GEN_10426 : _GEN_10374; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10459 = _T_1600 ? _GEN_10427 : _GEN_10375; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 118:26]
  wire [63:0] _GEN_10460 = csrAddr == 12'h301 ? _T_1802 : _GEN_10376; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  next_csr_mstatus_mstatusOld_3_pad4 = _T_1802[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_sie = _T_1802[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_pad3 = _T_1802[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_mie = _T_1802[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_pad2 = _T_1802[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_spie = _T_1802[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_ube = _T_1802[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_mpie = _T_1802[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_spp = _T_1802[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_3_vs = _T_1802[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_3_mpp = _T_1802[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_3_fs = _T_1802[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_3_xs = _T_1802[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_mprv = _T_1802[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_sum = _T_1802[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_mxr = _T_1802[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_tvm = _T_1802[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_tw = _T_1802[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_tsr = _T_1802[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [8:0] next_csr_mstatus_mstatusOld_3_pad0 = _T_1802[31:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_3_uxl = _T_1802[33:32]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_3_sxl = _T_1802[35:34]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_sbe = _T_1802[36]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_mbe = _T_1802[37]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [24:0] next_csr_mstatus_mstatusOld_3_pad1 = _T_1802[62:38]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_3_sd = _T_1802[63]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [5:0] next_csr_mstatus_mstatusNew_lo_lo_3 = {next_csr_mstatus_mstatusOld_3_spie,
    next_csr_mstatus_mstatusOld_3_pad2,next_csr_mstatus_mstatusOld_3_mie,next_csr_mstatus_mstatusOld_3_pad3,
    next_csr_mstatus_mstatusOld_3_sie,next_csr_mstatus_mstatusOld_3_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [16:0] next_csr_mstatus_mstatusNew_lo_3 = {next_csr_mstatus_mstatusOld_3_xs,next_csr_mstatus_mstatusOld_3_fs,
    next_csr_mstatus_mstatusOld_3_mpp,next_csr_mstatus_mstatusOld_3_vs,next_csr_mstatus_mstatusOld_3_spp,
    next_csr_mstatus_mstatusOld_3_mpie,next_csr_mstatus_mstatusOld_3_ube,next_csr_mstatus_mstatusNew_lo_lo_3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [5:0] next_csr_mstatus_mstatusNew_hi_lo_3 = {next_csr_mstatus_mstatusOld_3_tsr,next_csr_mstatus_mstatusOld_3_tw,
    next_csr_mstatus_mstatusOld_3_tvm,next_csr_mstatus_mstatusOld_3_mxr,next_csr_mstatus_mstatusOld_3_sum,
    next_csr_mstatus_mstatusOld_3_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [63:0] _next_csr_mstatus_mstatusNew_T_10 = {next_csr_mstatus_mstatusOld_3_sd,next_csr_mstatus_mstatusOld_3_pad1,
    next_csr_mstatus_mstatusOld_3_mbe,next_csr_mstatus_mstatusOld_3_sbe,next_csr_mstatus_mstatusOld_3_sxl,
    next_csr_mstatus_mstatusOld_3_uxl,next_csr_mstatus_mstatusOld_3_pad0,next_csr_mstatus_mstatusNew_hi_lo_3,
    next_csr_mstatus_mstatusNew_lo_3}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [63:0] next_csr_mstatus_mstatusNew_3 = {next_csr_mstatus_mstatusOld_3_fs == 2'h3,
    _next_csr_mstatus_mstatusNew_T_10[62:0]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:27]
  wire [63:0] _GEN_10461 = csrAddr == 12'h300 ? next_csr_mstatus_mstatusNew_3 : _GEN_10377; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10462 = csrAddr == 12'h340 ? _T_1802 : _GEN_10378; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10463 = csrAddr == 12'h305 ? _T_1802 : _GEN_10379; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10464 = csrAddr == 12'h306 ? _T_1802 : _GEN_10380; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _next_csr_mip_T_14 = _T_1802 & 64'h77f; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:80]
  wire [63:0] _next_csr_mip_T_15 = _next_csr_mip_T_1 | _next_csr_mip_T_14; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:72]
  wire [63:0] _GEN_10465 = csrAddr == 12'h344 ? _next_csr_mip_T_15 : _GEN_10381; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10466 = csrAddr == 12'h304 ? _T_1802 : _GEN_10382; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10468 = csrAddr == 12'h342 ? _T_1802 : _GEN_10384; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10469 = csrAddr == 12'h343 ? _T_1802 : _GEN_10385; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10470 = has_15 ? _GEN_10460 : _GEN_10376; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10471 = has_15 ? _GEN_10461 : _GEN_10377; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10472 = has_15 ? _GEN_10462 : _GEN_10378; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10473 = has_15 ? _GEN_10463 : _GEN_10379; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10474 = has_15 ? _GEN_10464 : _GEN_10380; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10475 = has_15 ? _GEN_10465 : _GEN_10381; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10476 = has_15 ? _GEN_10466 : _GEN_10382; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10478 = has_15 ? _GEN_10468 : _GEN_10384; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10479 = has_15 ? _GEN_10469 : _GEN_10385; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10483 = _T_1793 ? _GEN_10429 : _GEN_10345; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10484 = _T_1793 ? _GEN_10430 : _GEN_10346; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10485 = _T_1793 ? _GEN_10431 : _GEN_10347; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10486 = _T_1793 ? _GEN_10432 : _GEN_10348; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10487 = _T_1793 ? _GEN_10433 : _GEN_10349; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10488 = _T_1793 ? _GEN_10434 : _GEN_10350; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10489 = _T_1793 ? _GEN_10435 : _GEN_10351; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10490 = _T_1793 ? _GEN_10436 : _GEN_10352; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10491 = _T_1793 ? _GEN_10437 : _GEN_10353; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10492 = _T_1793 ? _GEN_10438 : _GEN_10354; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10493 = _T_1793 ? _GEN_10439 : _GEN_10355; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10494 = _T_1793 ? _GEN_10440 : _GEN_10356; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10495 = _T_1793 ? _GEN_10441 : _GEN_10357; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10496 = _T_1793 ? _GEN_10442 : _GEN_10358; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10497 = _T_1793 ? _GEN_10443 : _GEN_10359; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10498 = _T_1793 ? _GEN_10444 : _GEN_10360; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10499 = _T_1793 ? _GEN_10445 : _GEN_10361; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10500 = _T_1793 ? _GEN_10446 : _GEN_10362; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10501 = _T_1793 ? _GEN_10447 : _GEN_10363; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10502 = _T_1793 ? _GEN_10448 : _GEN_10364; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10503 = _T_1793 ? _GEN_10449 : _GEN_10365; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10504 = _T_1793 ? _GEN_10450 : _GEN_10366; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10505 = _T_1793 ? _GEN_10451 : _GEN_10367; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10506 = _T_1793 ? _GEN_10452 : _GEN_10368; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10507 = _T_1793 ? _GEN_10453 : _GEN_10369; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10508 = _T_1793 ? _GEN_10454 : _GEN_10370; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10509 = _T_1793 ? _GEN_10455 : _GEN_10371; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10510 = _T_1793 ? _GEN_10456 : _GEN_10372; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10511 = _T_1793 ? _GEN_10457 : _GEN_10373; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10512 = _T_1793 ? _GEN_10458 : _GEN_10374; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10513 = _T_1793 ? _GEN_10459 : _GEN_10375; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10514 = _T_1793 ? _GEN_10470 : _GEN_10376; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10515 = _T_1793 ? _GEN_10471 : _GEN_10377; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10516 = _T_1793 ? _GEN_10472 : _GEN_10378; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10517 = _T_1793 ? _GEN_10473 : _GEN_10379; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10518 = _T_1793 ? _GEN_10474 : _GEN_10380; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10519 = _T_1793 ? _GEN_10475 : _GEN_10381; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10520 = _T_1793 ? _GEN_10476 : _GEN_10382; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10522 = _T_1793 ? _GEN_10478 : _GEN_10384; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10523 = _T_1793 ? _GEN_10479 : _GEN_10385; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 117:27]
  wire [63:0] _GEN_10537 = _T_1709 ? _GEN_10483 : _GEN_10345; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10538 = _T_1709 ? _GEN_10484 : _GEN_10346; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10539 = _T_1709 ? _GEN_10485 : _GEN_10347; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10540 = _T_1709 ? _GEN_10486 : _GEN_10348; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10541 = _T_1709 ? _GEN_10487 : _GEN_10349; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10542 = _T_1709 ? _GEN_10488 : _GEN_10350; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10543 = _T_1709 ? _GEN_10489 : _GEN_10351; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10544 = _T_1709 ? _GEN_10490 : _GEN_10352; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10545 = _T_1709 ? _GEN_10491 : _GEN_10353; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10546 = _T_1709 ? _GEN_10492 : _GEN_10354; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10547 = _T_1709 ? _GEN_10493 : _GEN_10355; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10548 = _T_1709 ? _GEN_10494 : _GEN_10356; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10549 = _T_1709 ? _GEN_10495 : _GEN_10357; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10550 = _T_1709 ? _GEN_10496 : _GEN_10358; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10551 = _T_1709 ? _GEN_10497 : _GEN_10359; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10552 = _T_1709 ? _GEN_10498 : _GEN_10360; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10553 = _T_1709 ? _GEN_10499 : _GEN_10361; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10554 = _T_1709 ? _GEN_10500 : _GEN_10362; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10555 = _T_1709 ? _GEN_10501 : _GEN_10363; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10556 = _T_1709 ? _GEN_10502 : _GEN_10364; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10557 = _T_1709 ? _GEN_10503 : _GEN_10365; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10558 = _T_1709 ? _GEN_10504 : _GEN_10366; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10559 = _T_1709 ? _GEN_10505 : _GEN_10367; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10560 = _T_1709 ? _GEN_10506 : _GEN_10368; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10561 = _T_1709 ? _GEN_10507 : _GEN_10369; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10562 = _T_1709 ? _GEN_10508 : _GEN_10370; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10563 = _T_1709 ? _GEN_10509 : _GEN_10371; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10564 = _T_1709 ? _GEN_10510 : _GEN_10372; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10565 = _T_1709 ? _GEN_10511 : _GEN_10373; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10566 = _T_1709 ? _GEN_10512 : _GEN_10374; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10567 = _T_1709 ? _GEN_10513 : _GEN_10375; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10568 = _T_1709 ? _GEN_10514 : _GEN_10376; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10569 = _T_1709 ? _GEN_10515 : _GEN_10377; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10570 = _T_1709 ? _GEN_10516 : _GEN_10378; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10571 = _T_1709 ? _GEN_10517 : _GEN_10379; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10572 = _T_1709 ? _GEN_10518 : _GEN_10380; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10573 = _T_1709 ? _GEN_10519 : _GEN_10381; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10574 = _T_1709 ? _GEN_10520 : _GEN_10382; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10576 = _T_1709 ? _GEN_10522 : _GEN_10384; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10577 = _T_1709 ? _GEN_10523 : _GEN_10385; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 114:24]
  wire [63:0] _GEN_10589 = 5'h1 == rd ? rData_3 : _GEN_10537; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10590 = 5'h2 == rd ? rData_3 : _GEN_10538; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10591 = 5'h3 == rd ? rData_3 : _GEN_10539; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10592 = 5'h4 == rd ? rData_3 : _GEN_10540; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10593 = 5'h5 == rd ? rData_3 : _GEN_10541; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10594 = 5'h6 == rd ? rData_3 : _GEN_10542; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10595 = 5'h7 == rd ? rData_3 : _GEN_10543; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10596 = 5'h8 == rd ? rData_3 : _GEN_10544; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10597 = 5'h9 == rd ? rData_3 : _GEN_10545; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10598 = 5'ha == rd ? rData_3 : _GEN_10546; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10599 = 5'hb == rd ? rData_3 : _GEN_10547; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10600 = 5'hc == rd ? rData_3 : _GEN_10548; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10601 = 5'hd == rd ? rData_3 : _GEN_10549; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10602 = 5'he == rd ? rData_3 : _GEN_10550; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10603 = 5'hf == rd ? rData_3 : _GEN_10551; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10604 = 5'h10 == rd ? rData_3 : _GEN_10552; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10605 = 5'h11 == rd ? rData_3 : _GEN_10553; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10606 = 5'h12 == rd ? rData_3 : _GEN_10554; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10607 = 5'h13 == rd ? rData_3 : _GEN_10555; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10608 = 5'h14 == rd ? rData_3 : _GEN_10556; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10609 = 5'h15 == rd ? rData_3 : _GEN_10557; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10610 = 5'h16 == rd ? rData_3 : _GEN_10558; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10611 = 5'h17 == rd ? rData_3 : _GEN_10559; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10612 = 5'h18 == rd ? rData_3 : _GEN_10560; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10613 = 5'h19 == rd ? rData_3 : _GEN_10561; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10614 = 5'h1a == rd ? rData_3 : _GEN_10562; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10615 = 5'h1b == rd ? rData_3 : _GEN_10563; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10616 = 5'h1c == rd ? rData_3 : _GEN_10564; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10617 = 5'h1d == rd ? rData_3 : _GEN_10565; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10618 = 5'h1e == rd ? rData_3 : _GEN_10566; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10619 = 5'h1f == rd ? rData_3 : _GEN_10567; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 128:{22,22}]
  wire [63:0] _GEN_10628 = csrAddr == 12'h301 ? _T_1761 : _GEN_10568; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  next_csr_mstatus_mstatusOld_4_pad4 = _T_1761[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_sie = _T_1761[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_pad3 = _T_1761[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_mie = _T_1761[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_pad2 = _T_1761[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_spie = _T_1761[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_ube = _T_1761[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_mpie = _T_1761[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_spp = _T_1761[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_4_vs = _T_1761[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_4_mpp = _T_1761[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_4_fs = _T_1761[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_4_xs = _T_1761[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_mprv = _T_1761[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_sum = _T_1761[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_mxr = _T_1761[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_tvm = _T_1761[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_tw = _T_1761[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_tsr = _T_1761[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [8:0] next_csr_mstatus_mstatusOld_4_pad0 = _T_1761[31:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_4_uxl = _T_1761[33:32]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_4_sxl = _T_1761[35:34]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_sbe = _T_1761[36]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_mbe = _T_1761[37]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [24:0] next_csr_mstatus_mstatusOld_4_pad1 = _T_1761[62:38]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_4_sd = _T_1761[63]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [5:0] next_csr_mstatus_mstatusNew_lo_lo_4 = {next_csr_mstatus_mstatusOld_4_spie,
    next_csr_mstatus_mstatusOld_4_pad2,next_csr_mstatus_mstatusOld_4_mie,next_csr_mstatus_mstatusOld_4_pad3,
    next_csr_mstatus_mstatusOld_4_sie,next_csr_mstatus_mstatusOld_4_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [16:0] next_csr_mstatus_mstatusNew_lo_4 = {next_csr_mstatus_mstatusOld_4_xs,next_csr_mstatus_mstatusOld_4_fs,
    next_csr_mstatus_mstatusOld_4_mpp,next_csr_mstatus_mstatusOld_4_vs,next_csr_mstatus_mstatusOld_4_spp,
    next_csr_mstatus_mstatusOld_4_mpie,next_csr_mstatus_mstatusOld_4_ube,next_csr_mstatus_mstatusNew_lo_lo_4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [5:0] next_csr_mstatus_mstatusNew_hi_lo_4 = {next_csr_mstatus_mstatusOld_4_tsr,next_csr_mstatus_mstatusOld_4_tw,
    next_csr_mstatus_mstatusOld_4_tvm,next_csr_mstatus_mstatusOld_4_mxr,next_csr_mstatus_mstatusOld_4_sum,
    next_csr_mstatus_mstatusOld_4_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [63:0] _next_csr_mstatus_mstatusNew_T_13 = {next_csr_mstatus_mstatusOld_4_sd,next_csr_mstatus_mstatusOld_4_pad1,
    next_csr_mstatus_mstatusOld_4_mbe,next_csr_mstatus_mstatusOld_4_sbe,next_csr_mstatus_mstatusOld_4_sxl,
    next_csr_mstatus_mstatusOld_4_uxl,next_csr_mstatus_mstatusOld_4_pad0,next_csr_mstatus_mstatusNew_hi_lo_4,
    next_csr_mstatus_mstatusNew_lo_4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [63:0] next_csr_mstatus_mstatusNew_4 = {next_csr_mstatus_mstatusOld_4_fs == 2'h3,
    _next_csr_mstatus_mstatusNew_T_13[62:0]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:27]
  wire [63:0] _GEN_10629 = csrAddr == 12'h300 ? next_csr_mstatus_mstatusNew_4 : _GEN_10569; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10630 = csrAddr == 12'h340 ? _T_1761 : _GEN_10570; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10631 = csrAddr == 12'h305 ? _T_1761 : _GEN_10571; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10632 = csrAddr == 12'h306 ? _T_1761 : _GEN_10572; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _next_csr_mip_T_18 = _T_1761 & 64'h77f; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:80]
  wire [63:0] _next_csr_mip_T_19 = _next_csr_mip_T_1 | _next_csr_mip_T_18; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:72]
  wire [63:0] _GEN_10633 = csrAddr == 12'h344 ? _next_csr_mip_T_19 : _GEN_10573; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10634 = csrAddr == 12'h304 ? _T_1761 : _GEN_10574; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10636 = csrAddr == 12'h342 ? _T_1761 : _GEN_10576; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10637 = csrAddr == 12'h343 ? _T_1761 : _GEN_10577; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10638 = has_15 ? _GEN_10628 : _GEN_10568; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10639 = has_15 ? _GEN_10629 : _GEN_10569; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10640 = has_15 ? _GEN_10630 : _GEN_10570; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10641 = has_15 ? _GEN_10631 : _GEN_10571; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10642 = has_15 ? _GEN_10632 : _GEN_10572; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10643 = has_15 ? _GEN_10633 : _GEN_10573; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10644 = has_15 ? _GEN_10634 : _GEN_10574; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10646 = has_15 ? _GEN_10636 : _GEN_10576; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10647 = has_15 ? _GEN_10637 : _GEN_10577; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10650 = _T_1794 ? _GEN_10638 : _GEN_10568; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [63:0] _GEN_10651 = _T_1794 ? _GEN_10639 : _GEN_10569; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [63:0] _GEN_10652 = _T_1794 ? _GEN_10640 : _GEN_10570; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [63:0] _GEN_10653 = _T_1794 ? _GEN_10641 : _GEN_10571; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [63:0] _GEN_10654 = _T_1794 ? _GEN_10642 : _GEN_10572; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [63:0] _GEN_10655 = _T_1794 ? _GEN_10643 : _GEN_10573; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [63:0] _GEN_10656 = _T_1794 ? _GEN_10644 : _GEN_10574; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [63:0] _GEN_10658 = _T_1794 ? _GEN_10646 : _GEN_10576; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [63:0] _GEN_10659 = _T_1794 ? _GEN_10647 : _GEN_10577; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 130:27]
  wire [63:0] _GEN_10663 = ~isIllegalWrite_4 ? _GEN_10589 : _GEN_10537; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10664 = ~isIllegalWrite_4 ? _GEN_10590 : _GEN_10538; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10665 = ~isIllegalWrite_4 ? _GEN_10591 : _GEN_10539; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10666 = ~isIllegalWrite_4 ? _GEN_10592 : _GEN_10540; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10667 = ~isIllegalWrite_4 ? _GEN_10593 : _GEN_10541; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10668 = ~isIllegalWrite_4 ? _GEN_10594 : _GEN_10542; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10669 = ~isIllegalWrite_4 ? _GEN_10595 : _GEN_10543; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10670 = ~isIllegalWrite_4 ? _GEN_10596 : _GEN_10544; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10671 = ~isIllegalWrite_4 ? _GEN_10597 : _GEN_10545; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10672 = ~isIllegalWrite_4 ? _GEN_10598 : _GEN_10546; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10673 = ~isIllegalWrite_4 ? _GEN_10599 : _GEN_10547; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10674 = ~isIllegalWrite_4 ? _GEN_10600 : _GEN_10548; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10675 = ~isIllegalWrite_4 ? _GEN_10601 : _GEN_10549; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10676 = ~isIllegalWrite_4 ? _GEN_10602 : _GEN_10550; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10677 = ~isIllegalWrite_4 ? _GEN_10603 : _GEN_10551; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10678 = ~isIllegalWrite_4 ? _GEN_10604 : _GEN_10552; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10679 = ~isIllegalWrite_4 ? _GEN_10605 : _GEN_10553; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10680 = ~isIllegalWrite_4 ? _GEN_10606 : _GEN_10554; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10681 = ~isIllegalWrite_4 ? _GEN_10607 : _GEN_10555; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10682 = ~isIllegalWrite_4 ? _GEN_10608 : _GEN_10556; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10683 = ~isIllegalWrite_4 ? _GEN_10609 : _GEN_10557; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10684 = ~isIllegalWrite_4 ? _GEN_10610 : _GEN_10558; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10685 = ~isIllegalWrite_4 ? _GEN_10611 : _GEN_10559; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10686 = ~isIllegalWrite_4 ? _GEN_10612 : _GEN_10560; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10687 = ~isIllegalWrite_4 ? _GEN_10613 : _GEN_10561; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10688 = ~isIllegalWrite_4 ? _GEN_10614 : _GEN_10562; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10689 = ~isIllegalWrite_4 ? _GEN_10615 : _GEN_10563; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10690 = ~isIllegalWrite_4 ? _GEN_10616 : _GEN_10564; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10691 = ~isIllegalWrite_4 ? _GEN_10617 : _GEN_10565; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10692 = ~isIllegalWrite_4 ? _GEN_10618 : _GEN_10566; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10693 = ~isIllegalWrite_4 ? _GEN_10619 : _GEN_10567; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10694 = ~isIllegalWrite_4 ? _GEN_10650 : _GEN_10568; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10695 = ~isIllegalWrite_4 ? _GEN_10651 : _GEN_10569; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10696 = ~isIllegalWrite_4 ? _GEN_10652 : _GEN_10570; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10697 = ~isIllegalWrite_4 ? _GEN_10653 : _GEN_10571; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10698 = ~isIllegalWrite_4 ? _GEN_10654 : _GEN_10572; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10699 = ~isIllegalWrite_4 ? _GEN_10655 : _GEN_10573; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10700 = ~isIllegalWrite_4 ? _GEN_10656 : _GEN_10574; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10702 = ~isIllegalWrite_4 ? _GEN_10658 : _GEN_10576; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10703 = ~isIllegalWrite_4 ? _GEN_10659 : _GEN_10577; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 127:49]
  wire [63:0] _GEN_10717 = _T_1743 ? _GEN_10663 : _GEN_10537; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10718 = _T_1743 ? _GEN_10664 : _GEN_10538; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10719 = _T_1743 ? _GEN_10665 : _GEN_10539; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10720 = _T_1743 ? _GEN_10666 : _GEN_10540; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10721 = _T_1743 ? _GEN_10667 : _GEN_10541; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10722 = _T_1743 ? _GEN_10668 : _GEN_10542; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10723 = _T_1743 ? _GEN_10669 : _GEN_10543; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10724 = _T_1743 ? _GEN_10670 : _GEN_10544; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10725 = _T_1743 ? _GEN_10671 : _GEN_10545; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10726 = _T_1743 ? _GEN_10672 : _GEN_10546; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10727 = _T_1743 ? _GEN_10673 : _GEN_10547; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10728 = _T_1743 ? _GEN_10674 : _GEN_10548; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10729 = _T_1743 ? _GEN_10675 : _GEN_10549; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10730 = _T_1743 ? _GEN_10676 : _GEN_10550; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10731 = _T_1743 ? _GEN_10677 : _GEN_10551; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10732 = _T_1743 ? _GEN_10678 : _GEN_10552; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10733 = _T_1743 ? _GEN_10679 : _GEN_10553; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10734 = _T_1743 ? _GEN_10680 : _GEN_10554; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10735 = _T_1743 ? _GEN_10681 : _GEN_10555; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10736 = _T_1743 ? _GEN_10682 : _GEN_10556; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10737 = _T_1743 ? _GEN_10683 : _GEN_10557; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10738 = _T_1743 ? _GEN_10684 : _GEN_10558; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10739 = _T_1743 ? _GEN_10685 : _GEN_10559; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10740 = _T_1743 ? _GEN_10686 : _GEN_10560; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10741 = _T_1743 ? _GEN_10687 : _GEN_10561; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10742 = _T_1743 ? _GEN_10688 : _GEN_10562; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10743 = _T_1743 ? _GEN_10689 : _GEN_10563; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10744 = _T_1743 ? _GEN_10690 : _GEN_10564; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10745 = _T_1743 ? _GEN_10691 : _GEN_10565; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10746 = _T_1743 ? _GEN_10692 : _GEN_10566; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10747 = _T_1743 ? _GEN_10693 : _GEN_10567; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10748 = _T_1743 ? _GEN_10694 : _GEN_10568; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10749 = _T_1743 ? _GEN_10695 : _GEN_10569; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10750 = _T_1743 ? _GEN_10696 : _GEN_10570; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10751 = _T_1743 ? _GEN_10697 : _GEN_10571; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10752 = _T_1743 ? _GEN_10698 : _GEN_10572; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10753 = _T_1743 ? _GEN_10699 : _GEN_10573; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10754 = _T_1743 ? _GEN_10700 : _GEN_10574; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10756 = _T_1743 ? _GEN_10702 : _GEN_10576; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10757 = _T_1743 ? _GEN_10703 : _GEN_10577; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 124:24]
  wire [63:0] _GEN_10769 = 5'h1 == rd ? rData_3 : _GEN_10717; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10770 = 5'h2 == rd ? rData_3 : _GEN_10718; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10771 = 5'h3 == rd ? rData_3 : _GEN_10719; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10772 = 5'h4 == rd ? rData_3 : _GEN_10720; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10773 = 5'h5 == rd ? rData_3 : _GEN_10721; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10774 = 5'h6 == rd ? rData_3 : _GEN_10722; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10775 = 5'h7 == rd ? rData_3 : _GEN_10723; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10776 = 5'h8 == rd ? rData_3 : _GEN_10724; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10777 = 5'h9 == rd ? rData_3 : _GEN_10725; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10778 = 5'ha == rd ? rData_3 : _GEN_10726; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10779 = 5'hb == rd ? rData_3 : _GEN_10727; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10780 = 5'hc == rd ? rData_3 : _GEN_10728; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10781 = 5'hd == rd ? rData_3 : _GEN_10729; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10782 = 5'he == rd ? rData_3 : _GEN_10730; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10783 = 5'hf == rd ? rData_3 : _GEN_10731; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10784 = 5'h10 == rd ? rData_3 : _GEN_10732; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10785 = 5'h11 == rd ? rData_3 : _GEN_10733; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10786 = 5'h12 == rd ? rData_3 : _GEN_10734; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10787 = 5'h13 == rd ? rData_3 : _GEN_10735; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10788 = 5'h14 == rd ? rData_3 : _GEN_10736; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10789 = 5'h15 == rd ? rData_3 : _GEN_10737; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10790 = 5'h16 == rd ? rData_3 : _GEN_10738; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10791 = 5'h17 == rd ? rData_3 : _GEN_10739; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10792 = 5'h18 == rd ? rData_3 : _GEN_10740; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10793 = 5'h19 == rd ? rData_3 : _GEN_10741; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10794 = 5'h1a == rd ? rData_3 : _GEN_10742; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10795 = 5'h1b == rd ? rData_3 : _GEN_10743; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10796 = 5'h1c == rd ? rData_3 : _GEN_10744; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10797 = 5'h1d == rd ? rData_3 : _GEN_10745; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10798 = 5'h1e == rd ? rData_3 : _GEN_10746; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10799 = 5'h1f == rd ? rData_3 : _GEN_10747; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 139:{22,22}]
  wire [63:0] _GEN_10808 = csrAddr == 12'h301 ? _T_1804 : _GEN_10748; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire  next_csr_mstatus_mstatusOld_5_pad4 = _T_1804[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_sie = _T_1804[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_pad3 = _T_1804[2]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_mie = _T_1804[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_pad2 = _T_1804[4]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_spie = _T_1804[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_ube = _T_1804[6]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_mpie = _T_1804[7]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_spp = _T_1804[8]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_5_vs = _T_1804[10:9]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_5_mpp = _T_1804[12:11]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_5_fs = _T_1804[14:13]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_5_xs = _T_1804[16:15]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_mprv = _T_1804[17]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_sum = _T_1804[18]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_mxr = _T_1804[19]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_tvm = _T_1804[20]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_tw = _T_1804[21]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_tsr = _T_1804[22]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [8:0] next_csr_mstatus_mstatusOld_5_pad0 = _T_1804[31:23]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_5_uxl = _T_1804[33:32]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [1:0] next_csr_mstatus_mstatusOld_5_sxl = _T_1804[35:34]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_sbe = _T_1804[36]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_mbe = _T_1804[37]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [24:0] next_csr_mstatus_mstatusOld_5_pad1 = _T_1804[62:38]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire  next_csr_mstatus_mstatusOld_5_sd = _T_1804[63]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 52:49]
  wire [5:0] next_csr_mstatus_mstatusNew_lo_lo_5 = {next_csr_mstatus_mstatusOld_5_spie,
    next_csr_mstatus_mstatusOld_5_pad2,next_csr_mstatus_mstatusOld_5_mie,next_csr_mstatus_mstatusOld_5_pad3,
    next_csr_mstatus_mstatusOld_5_sie,next_csr_mstatus_mstatusOld_5_pad4}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [16:0] next_csr_mstatus_mstatusNew_lo_5 = {next_csr_mstatus_mstatusOld_5_xs,next_csr_mstatus_mstatusOld_5_fs,
    next_csr_mstatus_mstatusOld_5_mpp,next_csr_mstatus_mstatusOld_5_vs,next_csr_mstatus_mstatusOld_5_spp,
    next_csr_mstatus_mstatusOld_5_mpie,next_csr_mstatus_mstatusOld_5_ube,next_csr_mstatus_mstatusNew_lo_lo_5}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [5:0] next_csr_mstatus_mstatusNew_hi_lo_5 = {next_csr_mstatus_mstatusOld_5_tsr,next_csr_mstatus_mstatusOld_5_tw,
    next_csr_mstatus_mstatusOld_5_tvm,next_csr_mstatus_mstatusOld_5_mxr,next_csr_mstatus_mstatusOld_5_sum,
    next_csr_mstatus_mstatusOld_5_mprv}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [63:0] _next_csr_mstatus_mstatusNew_T_16 = {next_csr_mstatus_mstatusOld_5_sd,next_csr_mstatus_mstatusOld_5_pad1,
    next_csr_mstatus_mstatusOld_5_mbe,next_csr_mstatus_mstatusOld_5_sbe,next_csr_mstatus_mstatusOld_5_sxl,
    next_csr_mstatus_mstatusOld_5_uxl,next_csr_mstatus_mstatusOld_5_pad0,next_csr_mstatus_mstatusNew_hi_lo_5,
    next_csr_mstatus_mstatusNew_lo_5}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:66]
  wire [63:0] next_csr_mstatus_mstatusNew_5 = {next_csr_mstatus_mstatusOld_5_fs == 2'h3,
    _next_csr_mstatus_mstatusNew_T_16[62:0]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSR.scala 65:27]
  wire [63:0] _GEN_10809 = csrAddr == 12'h300 ? next_csr_mstatus_mstatusNew_5 : _GEN_10749; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10810 = csrAddr == 12'h340 ? _T_1804 : _GEN_10750; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10811 = csrAddr == 12'h305 ? _T_1804 : _GEN_10751; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10812 = csrAddr == 12'h306 ? _T_1804 : _GEN_10752; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _next_csr_mip_T_22 = _T_1804 & 64'h77f; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:80]
  wire [63:0] _next_csr_mip_T_23 = _next_csr_mip_T_1 | _next_csr_mip_T_22; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 70:72]
  wire [63:0] _GEN_10813 = csrAddr == 12'h344 ? _next_csr_mip_T_23 : _GEN_10753; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10814 = csrAddr == 12'h304 ? _T_1804 : _GEN_10754; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10816 = csrAddr == 12'h342 ? _T_1804 : _GEN_10756; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10817 = csrAddr == 12'h343 ? _T_1804 : _GEN_10757; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 67:34 70:21]
  wire [63:0] _GEN_10818 = has_15 ? _GEN_10808 : _GEN_10748; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10819 = has_15 ? _GEN_10809 : _GEN_10749; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10820 = has_15 ? _GEN_10810 : _GEN_10750; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10821 = has_15 ? _GEN_10811 : _GEN_10751; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10822 = has_15 ? _GEN_10812 : _GEN_10752; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10823 = has_15 ? _GEN_10813 : _GEN_10753; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10824 = has_15 ? _GEN_10814 : _GEN_10754; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10826 = has_15 ? _GEN_10816 : _GEN_10756; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10827 = has_15 ? _GEN_10817 : _GEN_10757; // @[src/main/scala/rvspeccore/core/spec/instset/csr/CSRSupport.scala 62:15]
  wire [63:0] _GEN_10830 = rs1 != 5'h0 ? _GEN_10818 : _GEN_10748; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [63:0] _GEN_10831 = rs1 != 5'h0 ? _GEN_10819 : _GEN_10749; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [63:0] _GEN_10832 = rs1 != 5'h0 ? _GEN_10820 : _GEN_10750; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [63:0] _GEN_10833 = rs1 != 5'h0 ? _GEN_10821 : _GEN_10751; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [63:0] _GEN_10834 = rs1 != 5'h0 ? _GEN_10822 : _GEN_10752; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [63:0] _GEN_10835 = rs1 != 5'h0 ? _GEN_10823 : _GEN_10753; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [63:0] _GEN_10836 = rs1 != 5'h0 ? _GEN_10824 : _GEN_10754; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [63:0] _GEN_10838 = rs1 != 5'h0 ? _GEN_10826 : _GEN_10756; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [63:0] _GEN_10839 = rs1 != 5'h0 ? _GEN_10827 : _GEN_10757; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 140:27]
  wire [63:0] _GEN_10843 = ~isIllegalWrite_5 ? _GEN_10769 : _GEN_10717; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10844 = ~isIllegalWrite_5 ? _GEN_10770 : _GEN_10718; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10845 = ~isIllegalWrite_5 ? _GEN_10771 : _GEN_10719; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10846 = ~isIllegalWrite_5 ? _GEN_10772 : _GEN_10720; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10847 = ~isIllegalWrite_5 ? _GEN_10773 : _GEN_10721; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10848 = ~isIllegalWrite_5 ? _GEN_10774 : _GEN_10722; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10849 = ~isIllegalWrite_5 ? _GEN_10775 : _GEN_10723; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10850 = ~isIllegalWrite_5 ? _GEN_10776 : _GEN_10724; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10851 = ~isIllegalWrite_5 ? _GEN_10777 : _GEN_10725; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10852 = ~isIllegalWrite_5 ? _GEN_10778 : _GEN_10726; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10853 = ~isIllegalWrite_5 ? _GEN_10779 : _GEN_10727; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10854 = ~isIllegalWrite_5 ? _GEN_10780 : _GEN_10728; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10855 = ~isIllegalWrite_5 ? _GEN_10781 : _GEN_10729; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10856 = ~isIllegalWrite_5 ? _GEN_10782 : _GEN_10730; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10857 = ~isIllegalWrite_5 ? _GEN_10783 : _GEN_10731; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10858 = ~isIllegalWrite_5 ? _GEN_10784 : _GEN_10732; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10859 = ~isIllegalWrite_5 ? _GEN_10785 : _GEN_10733; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10860 = ~isIllegalWrite_5 ? _GEN_10786 : _GEN_10734; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10861 = ~isIllegalWrite_5 ? _GEN_10787 : _GEN_10735; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10862 = ~isIllegalWrite_5 ? _GEN_10788 : _GEN_10736; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10863 = ~isIllegalWrite_5 ? _GEN_10789 : _GEN_10737; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10864 = ~isIllegalWrite_5 ? _GEN_10790 : _GEN_10738; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10865 = ~isIllegalWrite_5 ? _GEN_10791 : _GEN_10739; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10866 = ~isIllegalWrite_5 ? _GEN_10792 : _GEN_10740; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10867 = ~isIllegalWrite_5 ? _GEN_10793 : _GEN_10741; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10868 = ~isIllegalWrite_5 ? _GEN_10794 : _GEN_10742; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10869 = ~isIllegalWrite_5 ? _GEN_10795 : _GEN_10743; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10870 = ~isIllegalWrite_5 ? _GEN_10796 : _GEN_10744; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10871 = ~isIllegalWrite_5 ? _GEN_10797 : _GEN_10745; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10872 = ~isIllegalWrite_5 ? _GEN_10798 : _GEN_10746; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10873 = ~isIllegalWrite_5 ? _GEN_10799 : _GEN_10747; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10874 = ~isIllegalWrite_5 ? _GEN_10830 : _GEN_10748; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10875 = ~isIllegalWrite_5 ? _GEN_10831 : _GEN_10749; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10876 = ~isIllegalWrite_5 ? _GEN_10832 : _GEN_10750; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10877 = ~isIllegalWrite_5 ? _GEN_10833 : _GEN_10751; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10878 = ~isIllegalWrite_5 ? _GEN_10834 : _GEN_10752; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10879 = ~isIllegalWrite_5 ? _GEN_10835 : _GEN_10753; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10880 = ~isIllegalWrite_5 ? _GEN_10836 : _GEN_10754; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10882 = ~isIllegalWrite_5 ? _GEN_10838 : _GEN_10756; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10883 = ~isIllegalWrite_5 ? _GEN_10839 : _GEN_10757; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 138:27]
  wire [63:0] _GEN_10897 = _T_1786 ? _GEN_10843 : _GEN_10717; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10898 = _T_1786 ? _GEN_10844 : _GEN_10718; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10899 = _T_1786 ? _GEN_10845 : _GEN_10719; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10900 = _T_1786 ? _GEN_10846 : _GEN_10720; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10901 = _T_1786 ? _GEN_10847 : _GEN_10721; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10902 = _T_1786 ? _GEN_10848 : _GEN_10722; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10903 = _T_1786 ? _GEN_10849 : _GEN_10723; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10904 = _T_1786 ? _GEN_10850 : _GEN_10724; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10905 = _T_1786 ? _GEN_10851 : _GEN_10725; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10906 = _T_1786 ? _GEN_10852 : _GEN_10726; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10907 = _T_1786 ? _GEN_10853 : _GEN_10727; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10908 = _T_1786 ? _GEN_10854 : _GEN_10728; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10909 = _T_1786 ? _GEN_10855 : _GEN_10729; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10910 = _T_1786 ? _GEN_10856 : _GEN_10730; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10911 = _T_1786 ? _GEN_10857 : _GEN_10731; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10912 = _T_1786 ? _GEN_10858 : _GEN_10732; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10913 = _T_1786 ? _GEN_10859 : _GEN_10733; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10914 = _T_1786 ? _GEN_10860 : _GEN_10734; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10915 = _T_1786 ? _GEN_10861 : _GEN_10735; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10916 = _T_1786 ? _GEN_10862 : _GEN_10736; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10917 = _T_1786 ? _GEN_10863 : _GEN_10737; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10918 = _T_1786 ? _GEN_10864 : _GEN_10738; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10919 = _T_1786 ? _GEN_10865 : _GEN_10739; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10920 = _T_1786 ? _GEN_10866 : _GEN_10740; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10921 = _T_1786 ? _GEN_10867 : _GEN_10741; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10922 = _T_1786 ? _GEN_10868 : _GEN_10742; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10923 = _T_1786 ? _GEN_10869 : _GEN_10743; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10924 = _T_1786 ? _GEN_10870 : _GEN_10744; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10925 = _T_1786 ? _GEN_10871 : _GEN_10745; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10926 = _T_1786 ? _GEN_10872 : _GEN_10746; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10927 = _T_1786 ? _GEN_10873 : _GEN_10747; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10928 = _T_1786 ? _GEN_10874 : _GEN_10748; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10929 = _T_1786 ? _GEN_10875 : _GEN_10749; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10930 = _T_1786 ? _GEN_10876 : _GEN_10750; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10931 = _T_1786 ? _GEN_10877 : _GEN_10751; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10932 = _T_1786 ? _GEN_10878 : _GEN_10752; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10933 = _T_1786 ? _GEN_10879 : _GEN_10753; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10934 = _T_1786 ? _GEN_10880 : _GEN_10754; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10936 = _T_1786 ? _GEN_10882 : _GEN_10756; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire [63:0] _GEN_10937 = _T_1786 ? _GEN_10883 : _GEN_10757; // @[src/main/scala/rvspeccore/core/spec/instset/ZicsrExtension.scala 135:24]
  wire  _GEN_10950 = 2'h1 == io_now_csr_stvec[1:0] | _GEN_9816; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 316:29]
  wire  _GEN_10952 = 2'h0 == io_now_csr_stvec[1:0] | _GEN_10950; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 311:29]
  wire  _GEN_10975 = 8'h40 == io_now_csr_MXLEN ? _GEN_10952 : _GEN_9816; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire  _GEN_10985 = 8'h20 == io_now_csr_MXLEN ? _GEN_10952 : _GEN_10975; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire  _GEN_10993 = 2'h1 == io_now_csr_mtvec[1:0] | _GEN_9816; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 242:29]
  wire  _GEN_10995 = 2'h0 == io_now_csr_mtvec[1:0] | _GEN_10993; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 237:29]
  wire  _GEN_11015 = _T_1846 ? _GEN_10995 : _GEN_9816; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire  _GEN_11025 = _T_1829 ? _GEN_10995 : _GEN_11015; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire  _GEN_11036 = delegS ? _GEN_10985 : _GEN_11025; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire  _GEN_11053 = raiseExceptionIntr ? _GEN_11036 : _GEN_9816; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire  global_data_setpc = io_valid & _GEN_11053; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 113:21]
  wire [2:0] _next_pc_T_32 = inst[1:0] == 2'h3 ? 3'h4 : 3'h2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 154:32]
  wire [63:0] _GEN_11256 = {{61'd0}, _next_pc_T_32}; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 154:27]
  wire [63:0] _next_pc_T_34 = io_now_pc + _GEN_11256; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 154:27]
  wire [63:0] _GEN_10938 = ~global_data_setpc ? _next_pc_T_34 : _GEN_9817; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 150:30 154:17]
  wire [31:0] _next_csr_scause_T_1 = {1'h0,25'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 252:29]
  wire  mstatusNew_2_sie = delegS ? 1'h0 : io_now_csr_mstatus[1]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  mstatusNew_2_spie = delegS ? io_now_csr_mstatus[1] : io_now_csr_mstatus[5]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  mstatusNew_2_mie = delegS & io_now_csr_mstatus[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire [5:0] next_csr_mstatus_lo_lo_2 = {mstatusNew_2_spie,io_now_csr_mstatus[4],mstatusNew_2_mie,io_now_csr_mstatus[2],
    mstatusNew_2_sie,io_now_csr_mstatus[0]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [1:0] _GEN_11028 = delegS ? io_now_internal_privilegeMode : {{1'd0}, io_now_csr_mstatus[8]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire  mstatusNew_2_spp = _GEN_11028[0]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 159:30]
  wire  mstatusNew_2_mpie = delegS ? io_now_csr_mstatus[7] : io_now_csr_mstatus[3]; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire [1:0] mstatusNew_2_mpp = delegS ? next_reg_mstatusStruct_10_mpp : io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 159:30]
  wire [16:0] next_csr_mstatus_lo_2 = {io_now_csr_mstatus[16:15],io_now_csr_mstatus[14:13],mstatusNew_2_mpp,
    io_now_csr_mstatus[10:9],mstatusNew_2_spp,mstatusNew_2_mpie,io_now_csr_mstatus[6],next_csr_mstatus_lo_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire [63:0] _next_csr_mstatus_T_38 = {io_now_csr_mstatus[63],io_now_csr_mstatus[62:38],io_now_csr_mstatus[37],
    io_now_csr_mstatus[36],io_now_csr_mstatus[35:34],io_now_csr_mstatus[33:32],io_now_csr_mstatus[31:23],
    next_csr_mstatus_hi_lo_1,next_csr_mstatus_lo_2}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 260:49]
  wire  _T_1830 = 6'h2 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [31:0] _GEN_10941 = inst[1:0] != 2'h3 ? {{16'd0}, inst[15:0]} : inst; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 271:{45,62} 272:41]
  wire  _T_1833 = 6'h1 == exceptionNO; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29]
  wire [63:0] mem_read_addr = io_valid ? _GEN_8270 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [63:0] _GEN_10944 = 6'h4 == exceptionNO ? mem_read_addr : 64'h0; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29 296:26 259:35]
  wire [63:0] mem_write_addr = io_valid ? _GEN_8504 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  wire [63:0] _GEN_10945 = 6'h6 == exceptionNO ? mem_write_addr : _GEN_10944; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29 292:26]
  wire [63:0] _GEN_10946 = 6'hb == exceptionNO ? 64'h0 : _GEN_10945; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 263:29 288:26]
  wire [31:0] _next_pc_T_36 = {io_now_csr_stvec[31:2], 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 312:62]
  wire [31:0] _next_pc_T_38 = {26'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [31:0] _GEN_11257 = {{2'd0}, io_now_csr_stvec[31:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:60]
  wire [31:0] _next_pc_T_40 = _GEN_11257 + _next_pc_T_38; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:60]
  wire [33:0] _next_pc_T_41 = {_next_pc_T_40, 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:92]
  wire [63:0] _GEN_10951 = 2'h1 == io_now_csr_stvec[1:0] ? {{30'd0}, _next_pc_T_41} : _GEN_10938; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 317:29]
  wire [63:0] _GEN_10953 = 2'h0 == io_now_csr_stvec[1:0] ? {{32'd0}, _next_pc_T_36} : _GEN_10951; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 312:29]
  wire [63:0] _next_csr_scause_T_3 = {1'h0,57'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 252:29]
  wire [63:0] _next_pc_T_43 = {io_now_csr_stvec[63:2], 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 312:62]
  wire [63:0] _next_pc_T_45 = {58'h0,exceptionNO}; // @[src/main/scala/rvspeccore/core/tool/BitTool.scala 21:10]
  wire [63:0] _GEN_11258 = {{2'd0}, io_now_csr_stvec[63:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:60]
  wire [63:0] _next_pc_T_47 = _GEN_11258 + _next_pc_T_45; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:60]
  wire [65:0] _next_pc_T_48 = {_next_pc_T_47, 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 317:92]
  wire [65:0] _GEN_10964 = 2'h1 == io_now_csr_stvec[1:0] ? _next_pc_T_48 : {{2'd0}, _GEN_10938}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 317:29]
  wire [65:0] _GEN_10966 = 2'h0 == io_now_csr_stvec[1:0] ? {{2'd0}, _next_pc_T_43} : _GEN_10964; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 308:35 312:29]
  wire [63:0] _GEN_10967 = 8'h40 == io_now_csr_MXLEN ? _next_csr_scause_T_3 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 252:23]
  wire [65:0] _GEN_10976 = 8'h40 == io_now_csr_MXLEN ? _GEN_10966 : {{2'd0}, _GEN_10938}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire [63:0] _GEN_10977 = 8'h20 == io_now_csr_MXLEN ? {{32'd0}, _next_csr_scause_T_1} : _GEN_10967; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29 252:23]
  wire [65:0] _GEN_10986 = 8'h20 == io_now_csr_MXLEN ? {{2'd0}, _GEN_10953} : _GEN_10976; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 166:29]
  wire [63:0] _GEN_10991 = _T_1833 ? {{32'd0}, _GEN_10941} : _GEN_10946; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29]
  wire [63:0] _GEN_10992 = _T_1830 ? 64'h0 : _GEN_10991; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 196:29 199:26]
  wire [31:0] _next_pc_T_50 = {io_now_csr_mtvec[31:2], 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 238:62]
  wire [31:0] _GEN_11259 = {{2'd0}, io_now_csr_mtvec[31:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:60]
  wire [31:0] _next_pc_T_54 = _GEN_11259 + _next_pc_T_38; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:60]
  wire [33:0] _next_pc_T_55 = {_next_pc_T_54, 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:92]
  wire [63:0] _GEN_10994 = 2'h1 == io_now_csr_mtvec[1:0] ? {{30'd0}, _next_pc_T_55} : _GEN_10938; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 243:29]
  wire [63:0] _GEN_10996 = 2'h0 == io_now_csr_mtvec[1:0] ? {{32'd0}, _next_pc_T_50} : _GEN_10994; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 238:29]
  wire [63:0] _next_pc_T_57 = {io_now_csr_mtvec[63:2], 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 238:62]
  wire [63:0] _GEN_11260 = {{2'd0}, io_now_csr_mtvec[63:2]}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:60]
  wire [63:0] _next_pc_T_61 = _GEN_11260 + _next_pc_T_45; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:60]
  wire [65:0] _next_pc_T_62 = {_next_pc_T_61, 2'h0}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 243:92]
  wire [65:0] _GEN_11004 = 2'h1 == io_now_csr_mtvec[1:0] ? _next_pc_T_62 : {{2'd0}, _GEN_10938}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 243:29]
  wire [65:0] _GEN_11006 = 2'h0 == io_now_csr_mtvec[1:0] ? {{2'd0}, _next_pc_T_57} : _GEN_11004; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 234:35 238:29]
  wire [63:0] _GEN_11007 = _T_1846 ? _next_csr_scause_T_3 : _GEN_10936; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 185:35]
  wire [63:0] _GEN_11013 = _T_1846 ? _GEN_10992 : _GEN_10937; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire [65:0] _GEN_11016 = _T_1846 ? _GEN_11006 : {{2'd0}, _GEN_10938}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire [63:0] _GEN_11017 = _T_1829 ? {{32'd0}, _next_csr_scause_T_1} : _GEN_11007; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29 185:35]
  wire [63:0] _GEN_11023 = _T_1829 ? _GEN_10992 : _GEN_11013; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire [65:0] _GEN_11026 = _T_1829 ? {{2'd0}, _GEN_10996} : _GEN_11016; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 176:29]
  wire [63:0] _GEN_11032 = delegS ? _GEN_10977 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 src/main/scala/rvspeccore/core/RiscvCore.scala 111:21]
  wire [63:0] _GEN_11049 = raiseExceptionIntr ? _GEN_11032 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 111:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [63:0] next_csr_scause = io_valid ? _GEN_11049 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [63:0] _GEN_11041 = delegS ? _GEN_10936 : _GEN_11017; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [63:0] _GEN_11055 = raiseExceptionIntr ? _GEN_11041 : _GEN_10936; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [63:0] next_csr_mcause = io_valid ? _GEN_11055 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  wire [63:0] _GEN_11027 = delegS ? next_csr_scause : next_csr_mcause; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18 161:35 171:35]
  wire [1:0] _GEN_11031 = delegS ? 2'h1 : 2'h3; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [65:0] _GEN_11037 = delegS ? _GEN_10986 : _GEN_11026; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [63:0] _GEN_11043 = delegS ? _GEN_10937 : _GEN_11023; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 160:18]
  wire [63:0] _GEN_11045 = raiseExceptionIntr ? _GEN_11027 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [63:0] _GEN_11046 = raiseExceptionIntr ? io_now_pc : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30 151:25]
  wire [63:0] _GEN_11047 = raiseExceptionIntr ? {{32'd0}, inst} : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 114:21 src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30 152:25]
  wire [1:0] _GEN_11048 = raiseExceptionIntr ? _GEN_11031 : _GEN_9813; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [63:0] _GEN_11052 = raiseExceptionIntr ? _next_csr_mstatus_T_38 : _GEN_10929; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30 181:22]
  wire [65:0] _GEN_11054 = raiseExceptionIntr ? _GEN_11037 : {{2'd0}, _GEN_10938}; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [63:0] _GEN_11057 = raiseExceptionIntr ? _GEN_11043 : _GEN_10937; // @[src/main/scala/rvspeccore/core/spec/instset/csr/ExceptionSupport.scala 136:30]
  wire [65:0] _GEN_11119 = io_valid ? _GEN_11054 : {{2'd0}, io_now_pc}; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_mem_read_valid = io_valid & _GEN_8256; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_read_addr = io_valid ? _GEN_8270 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_read_memWidth = io_valid ? _GEN_8273 : 7'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_write_valid = io_valid & _GEN_8490; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_write_addr = io_valid ? _GEN_8504 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_write_memWidth = io_valid ? _GEN_8507 : 7'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_mem_write_data = io_valid ? _GEN_8508 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 119:7]
  assign io_tlb_Anotherread_0_valid = io_valid & _GEN_8491; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 123:18]
  assign io_tlb_Anotherread_0_addr = io_valid ? _GEN_8492 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 123:18]
  assign io_tlb_Anotherread_1_valid = io_valid & _GEN_8494; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 123:18]
  assign io_tlb_Anotherread_1_addr = io_valid ? _GEN_8495 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 123:18]
  assign io_tlb_Anotherread_2_valid = io_valid & _GEN_8497; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 123:18]
  assign io_tlb_Anotherread_2_addr = io_valid ? _GEN_8498 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 120:13 123:18]
  assign io_next_reg_0 = io_valid ? 64'h0 : io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 148:17 111:21]
  assign io_next_reg_1 = io_valid ? _GEN_10897 : io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_2 = io_valid ? _GEN_10898 : io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_3 = io_valid ? _GEN_10899 : io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_4 = io_valid ? _GEN_10900 : io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_5 = io_valid ? _GEN_10901 : io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_6 = io_valid ? _GEN_10902 : io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_7 = io_valid ? _GEN_10903 : io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_8 = io_valid ? _GEN_10904 : io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_9 = io_valid ? _GEN_10905 : io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_10 = io_valid ? _GEN_10906 : io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_11 = io_valid ? _GEN_10907 : io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_12 = io_valid ? _GEN_10908 : io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_13 = io_valid ? _GEN_10909 : io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_14 = io_valid ? _GEN_10910 : io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_15 = io_valid ? _GEN_10911 : io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_16 = io_valid ? _GEN_10912 : io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_17 = io_valid ? _GEN_10913 : io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_18 = io_valid ? _GEN_10914 : io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_19 = io_valid ? _GEN_10915 : io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_20 = io_valid ? _GEN_10916 : io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_21 = io_valid ? _GEN_10917 : io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_22 = io_valid ? _GEN_10918 : io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_23 = io_valid ? _GEN_10919 : io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_24 = io_valid ? _GEN_10920 : io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_25 = io_valid ? _GEN_10921 : io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_26 = io_valid ? _GEN_10922 : io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_27 = io_valid ? _GEN_10923 : io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_28 = io_valid ? _GEN_10924 : io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_29 = io_valid ? _GEN_10925 : io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_30 = io_valid ? _GEN_10926 : io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_reg_31 = io_valid ? _GEN_10927 : io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_pc = _GEN_11119[63:0]; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 18:18]
  assign io_next_csr_misa = io_valid ? _GEN_10928 : io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mvendorid = io_now_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_marchid = io_now_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mimpid = io_now_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mhartid = io_now_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mstatus = io_valid ? _GEN_11052 : io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mscratch = io_valid ? _GEN_10930 : io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mtvec = io_valid ? _GEN_10931 : io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mcounteren = io_valid ? _GEN_10932 : io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_medeleg = io_now_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_mip = io_valid ? _GEN_10933 : io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mie = io_valid ? _GEN_10934 : io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mepc = io_valid ? _GEN_11056 : io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mcause = io_valid ? _GEN_11055 : io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_mtval = io_valid ? _GEN_11057 : io_now_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_scause = io_valid ? _GEN_11049 : io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_stvec = io_now_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_sepc = io_valid ? _GEN_11050 : io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_next_csr_satp = io_now_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_MXLEN = io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_csr_IALIGN = io_now_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 17:18 109:7]
  assign io_next_internal_privilegeMode = io_valid ? _GEN_11048 : io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 111:21]
  assign io_event_valid = io_valid & raiseExceptionIntr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  assign io_event_cause = io_valid ? _GEN_11045 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  assign io_event_exceptionPC = io_valid ? _GEN_11046 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
  assign io_event_exceptionInst = io_valid ? _GEN_11047 : 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 123:18 114:21]
endmodule
module RiscvCore(
  input         clock,
  input         reset,
  input  [31:0] io_inst, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  input         io_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output        io_mem_read_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_mem_read_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [6:0]  io_mem_read_memWidth, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  input  [63:0] io_mem_read_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output        io_mem_write_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_mem_write_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [6:0]  io_mem_write_memWidth, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_mem_write_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output        io_tlb_Anotherread_0_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_tlb_Anotherread_0_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  input  [63:0] io_tlb_Anotherread_0_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output        io_tlb_Anotherread_1_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_tlb_Anotherread_1_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  input  [63:0] io_tlb_Anotherread_1_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output        io_tlb_Anotherread_2_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_tlb_Anotherread_2_addr, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  input  [63:0] io_tlb_Anotherread_2_data, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_now_pc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_0, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_1, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_2, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_3, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_4, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_5, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_6, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_7, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_8, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_9, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_10, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_11, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_12, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_13, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_14, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_15, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_16, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_17, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_18, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_19, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_20, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_21, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_22, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_23, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_24, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_25, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_26, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_27, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_28, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_29, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_30, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_reg_31, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_misa, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mvendorid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_marchid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mimpid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mhartid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mstatus, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mscratch, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mtvec, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mcounteren, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mip, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mie, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mepc, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mcause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_next_csr_mtval, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output        io_event_valid, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_event_cause, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_event_exceptionPC, // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
  output [63:0] io_event_exceptionInst // @[src/main/scala/rvspeccore/core/RiscvCore.scala 175:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] trans_io_inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_mem_read_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_mem_read_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [6:0] trans_io_mem_read_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_mem_read_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_mem_write_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_mem_write_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [6:0] trans_io_mem_write_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_mem_write_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_tlb_Anotherread_0_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_tlb_Anotherread_0_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_tlb_Anotherread_0_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_tlb_Anotherread_1_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_tlb_Anotherread_1_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_tlb_Anotherread_1_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_tlb_Anotherread_2_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_tlb_Anotherread_2_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_tlb_Anotherread_2_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_now_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_now_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_now_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [1:0] trans_io_now_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_next_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_next_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [7:0] trans_io_next_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [1:0] trans_io_next_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire  trans_io_event_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_event_cause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_event_exceptionPC; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  wire [63:0] trans_io_event_exceptionInst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
  reg [63:0] state_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [63:0] state_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [7:0] state_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [7:0] state_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  reg [1:0] state_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
  RiscvTrans trans ( // @[src/main/scala/rvspeccore/core/RiscvCore.scala 190:21]
    .io_inst(trans_io_inst),
    .io_valid(trans_io_valid),
    .io_mem_read_valid(trans_io_mem_read_valid),
    .io_mem_read_addr(trans_io_mem_read_addr),
    .io_mem_read_memWidth(trans_io_mem_read_memWidth),
    .io_mem_read_data(trans_io_mem_read_data),
    .io_mem_write_valid(trans_io_mem_write_valid),
    .io_mem_write_addr(trans_io_mem_write_addr),
    .io_mem_write_memWidth(trans_io_mem_write_memWidth),
    .io_mem_write_data(trans_io_mem_write_data),
    .io_tlb_Anotherread_0_valid(trans_io_tlb_Anotherread_0_valid),
    .io_tlb_Anotherread_0_addr(trans_io_tlb_Anotherread_0_addr),
    .io_tlb_Anotherread_0_data(trans_io_tlb_Anotherread_0_data),
    .io_tlb_Anotherread_1_valid(trans_io_tlb_Anotherread_1_valid),
    .io_tlb_Anotherread_1_addr(trans_io_tlb_Anotherread_1_addr),
    .io_tlb_Anotherread_1_data(trans_io_tlb_Anotherread_1_data),
    .io_tlb_Anotherread_2_valid(trans_io_tlb_Anotherread_2_valid),
    .io_tlb_Anotherread_2_addr(trans_io_tlb_Anotherread_2_addr),
    .io_tlb_Anotherread_2_data(trans_io_tlb_Anotherread_2_data),
    .io_now_reg_0(trans_io_now_reg_0),
    .io_now_reg_1(trans_io_now_reg_1),
    .io_now_reg_2(trans_io_now_reg_2),
    .io_now_reg_3(trans_io_now_reg_3),
    .io_now_reg_4(trans_io_now_reg_4),
    .io_now_reg_5(trans_io_now_reg_5),
    .io_now_reg_6(trans_io_now_reg_6),
    .io_now_reg_7(trans_io_now_reg_7),
    .io_now_reg_8(trans_io_now_reg_8),
    .io_now_reg_9(trans_io_now_reg_9),
    .io_now_reg_10(trans_io_now_reg_10),
    .io_now_reg_11(trans_io_now_reg_11),
    .io_now_reg_12(trans_io_now_reg_12),
    .io_now_reg_13(trans_io_now_reg_13),
    .io_now_reg_14(trans_io_now_reg_14),
    .io_now_reg_15(trans_io_now_reg_15),
    .io_now_reg_16(trans_io_now_reg_16),
    .io_now_reg_17(trans_io_now_reg_17),
    .io_now_reg_18(trans_io_now_reg_18),
    .io_now_reg_19(trans_io_now_reg_19),
    .io_now_reg_20(trans_io_now_reg_20),
    .io_now_reg_21(trans_io_now_reg_21),
    .io_now_reg_22(trans_io_now_reg_22),
    .io_now_reg_23(trans_io_now_reg_23),
    .io_now_reg_24(trans_io_now_reg_24),
    .io_now_reg_25(trans_io_now_reg_25),
    .io_now_reg_26(trans_io_now_reg_26),
    .io_now_reg_27(trans_io_now_reg_27),
    .io_now_reg_28(trans_io_now_reg_28),
    .io_now_reg_29(trans_io_now_reg_29),
    .io_now_reg_30(trans_io_now_reg_30),
    .io_now_reg_31(trans_io_now_reg_31),
    .io_now_pc(trans_io_now_pc),
    .io_now_csr_misa(trans_io_now_csr_misa),
    .io_now_csr_mvendorid(trans_io_now_csr_mvendorid),
    .io_now_csr_marchid(trans_io_now_csr_marchid),
    .io_now_csr_mimpid(trans_io_now_csr_mimpid),
    .io_now_csr_mhartid(trans_io_now_csr_mhartid),
    .io_now_csr_mstatus(trans_io_now_csr_mstatus),
    .io_now_csr_mscratch(trans_io_now_csr_mscratch),
    .io_now_csr_mtvec(trans_io_now_csr_mtvec),
    .io_now_csr_mcounteren(trans_io_now_csr_mcounteren),
    .io_now_csr_medeleg(trans_io_now_csr_medeleg),
    .io_now_csr_mip(trans_io_now_csr_mip),
    .io_now_csr_mie(trans_io_now_csr_mie),
    .io_now_csr_mepc(trans_io_now_csr_mepc),
    .io_now_csr_mcause(trans_io_now_csr_mcause),
    .io_now_csr_mtval(trans_io_now_csr_mtval),
    .io_now_csr_scause(trans_io_now_csr_scause),
    .io_now_csr_stvec(trans_io_now_csr_stvec),
    .io_now_csr_sepc(trans_io_now_csr_sepc),
    .io_now_csr_satp(trans_io_now_csr_satp),
    .io_now_csr_MXLEN(trans_io_now_csr_MXLEN),
    .io_now_csr_IALIGN(trans_io_now_csr_IALIGN),
    .io_now_internal_privilegeMode(trans_io_now_internal_privilegeMode),
    .io_next_reg_0(trans_io_next_reg_0),
    .io_next_reg_1(trans_io_next_reg_1),
    .io_next_reg_2(trans_io_next_reg_2),
    .io_next_reg_3(trans_io_next_reg_3),
    .io_next_reg_4(trans_io_next_reg_4),
    .io_next_reg_5(trans_io_next_reg_5),
    .io_next_reg_6(trans_io_next_reg_6),
    .io_next_reg_7(trans_io_next_reg_7),
    .io_next_reg_8(trans_io_next_reg_8),
    .io_next_reg_9(trans_io_next_reg_9),
    .io_next_reg_10(trans_io_next_reg_10),
    .io_next_reg_11(trans_io_next_reg_11),
    .io_next_reg_12(trans_io_next_reg_12),
    .io_next_reg_13(trans_io_next_reg_13),
    .io_next_reg_14(trans_io_next_reg_14),
    .io_next_reg_15(trans_io_next_reg_15),
    .io_next_reg_16(trans_io_next_reg_16),
    .io_next_reg_17(trans_io_next_reg_17),
    .io_next_reg_18(trans_io_next_reg_18),
    .io_next_reg_19(trans_io_next_reg_19),
    .io_next_reg_20(trans_io_next_reg_20),
    .io_next_reg_21(trans_io_next_reg_21),
    .io_next_reg_22(trans_io_next_reg_22),
    .io_next_reg_23(trans_io_next_reg_23),
    .io_next_reg_24(trans_io_next_reg_24),
    .io_next_reg_25(trans_io_next_reg_25),
    .io_next_reg_26(trans_io_next_reg_26),
    .io_next_reg_27(trans_io_next_reg_27),
    .io_next_reg_28(trans_io_next_reg_28),
    .io_next_reg_29(trans_io_next_reg_29),
    .io_next_reg_30(trans_io_next_reg_30),
    .io_next_reg_31(trans_io_next_reg_31),
    .io_next_pc(trans_io_next_pc),
    .io_next_csr_misa(trans_io_next_csr_misa),
    .io_next_csr_mvendorid(trans_io_next_csr_mvendorid),
    .io_next_csr_marchid(trans_io_next_csr_marchid),
    .io_next_csr_mimpid(trans_io_next_csr_mimpid),
    .io_next_csr_mhartid(trans_io_next_csr_mhartid),
    .io_next_csr_mstatus(trans_io_next_csr_mstatus),
    .io_next_csr_mscratch(trans_io_next_csr_mscratch),
    .io_next_csr_mtvec(trans_io_next_csr_mtvec),
    .io_next_csr_mcounteren(trans_io_next_csr_mcounteren),
    .io_next_csr_medeleg(trans_io_next_csr_medeleg),
    .io_next_csr_mip(trans_io_next_csr_mip),
    .io_next_csr_mie(trans_io_next_csr_mie),
    .io_next_csr_mepc(trans_io_next_csr_mepc),
    .io_next_csr_mcause(trans_io_next_csr_mcause),
    .io_next_csr_mtval(trans_io_next_csr_mtval),
    .io_next_csr_scause(trans_io_next_csr_scause),
    .io_next_csr_stvec(trans_io_next_csr_stvec),
    .io_next_csr_sepc(trans_io_next_csr_sepc),
    .io_next_csr_satp(trans_io_next_csr_satp),
    .io_next_csr_MXLEN(trans_io_next_csr_MXLEN),
    .io_next_csr_IALIGN(trans_io_next_csr_IALIGN),
    .io_next_internal_privilegeMode(trans_io_next_internal_privilegeMode),
    .io_event_valid(trans_io_event_valid),
    .io_event_cause(trans_io_event_cause),
    .io_event_exceptionPC(trans_io_event_exceptionPC),
    .io_event_exceptionInst(trans_io_event_exceptionInst)
  );
  assign io_mem_read_valid = trans_io_mem_read_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_read_addr = trans_io_mem_read_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_read_memWidth = trans_io_mem_read_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_write_valid = trans_io_mem_write_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_write_addr = trans_io_mem_write_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_write_memWidth = trans_io_mem_write_memWidth; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_mem_write_data = trans_io_mem_write_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign io_tlb_Anotherread_0_valid = trans_io_tlb_Anotherread_0_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 195:22]
  assign io_tlb_Anotherread_0_addr = trans_io_tlb_Anotherread_0_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 195:22]
  assign io_tlb_Anotherread_1_valid = trans_io_tlb_Anotherread_1_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 195:22]
  assign io_tlb_Anotherread_1_addr = trans_io_tlb_Anotherread_1_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 195:22]
  assign io_tlb_Anotherread_2_valid = trans_io_tlb_Anotherread_2_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 195:22]
  assign io_tlb_Anotherread_2_addr = trans_io_tlb_Anotherread_2_addr; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 195:22]
  assign io_now_pc = state_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 200:15]
  assign io_next_reg_0 = trans_io_next_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_1 = trans_io_next_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_2 = trans_io_next_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_3 = trans_io_next_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_4 = trans_io_next_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_5 = trans_io_next_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_6 = trans_io_next_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_7 = trans_io_next_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_8 = trans_io_next_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_9 = trans_io_next_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_10 = trans_io_next_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_11 = trans_io_next_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_12 = trans_io_next_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_13 = trans_io_next_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_14 = trans_io_next_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_15 = trans_io_next_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_16 = trans_io_next_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_17 = trans_io_next_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_18 = trans_io_next_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_19 = trans_io_next_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_20 = trans_io_next_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_21 = trans_io_next_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_22 = trans_io_next_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_23 = trans_io_next_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_24 = trans_io_next_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_25 = trans_io_next_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_26 = trans_io_next_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_27 = trans_io_next_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_28 = trans_io_next_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_29 = trans_io_next_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_30 = trans_io_next_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_reg_31 = trans_io_next_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_misa = trans_io_next_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mvendorid = trans_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_marchid = trans_io_next_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mimpid = trans_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mhartid = trans_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mstatus = trans_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mscratch = trans_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mtvec = trans_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mcounteren = trans_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mip = trans_io_next_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mie = trans_io_next_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mepc = trans_io_next_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mcause = trans_io_next_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_next_csr_mtval = trans_io_next_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 201:15]
  assign io_event_valid = trans_io_event_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign io_event_cause = trans_io_event_cause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign io_event_exceptionPC = trans_io_event_exceptionPC; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign io_event_exceptionInst = trans_io_event_exceptionInst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 202:15]
  assign trans_io_inst = io_inst; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 192:18]
  assign trans_io_valid = io_valid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 193:18]
  assign trans_io_mem_read_data = io_mem_read_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 194:16]
  assign trans_io_tlb_Anotherread_0_data = io_tlb_Anotherread_0_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 195:22]
  assign trans_io_tlb_Anotherread_1_data = io_tlb_Anotherread_1_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 195:22]
  assign trans_io_tlb_Anotherread_2_data = io_tlb_Anotherread_2_data; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 195:22]
  assign trans_io_now_reg_0 = state_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_1 = state_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_2 = state_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_3 = state_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_4 = state_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_5 = state_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_6 = state_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_7 = state_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_8 = state_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_9 = state_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_10 = state_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_11 = state_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_12 = state_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_13 = state_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_14 = state_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_15 = state_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_16 = state_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_17 = state_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_18 = state_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_19 = state_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_20 = state_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_21 = state_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_22 = state_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_23 = state_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_24 = state_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_25 = state_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_26 = state_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_27 = state_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_28 = state_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_29 = state_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_30 = state_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_reg_31 = state_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_pc = state_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_misa = state_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mvendorid = state_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_marchid = state_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mimpid = state_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mhartid = state_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mstatus = state_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mscratch = state_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mtvec = state_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mcounteren = state_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_medeleg = state_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mip = state_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mie = state_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mepc = state_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mcause = state_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_mtval = state_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_scause = state_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_stvec = state_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_sepc = state_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_satp = state_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_MXLEN = state_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_csr_IALIGN = state_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  assign trans_io_now_internal_privilegeMode = state_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 197:16]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_0 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_0 <= trans_io_next_reg_0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_1 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_1 <= trans_io_next_reg_1; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_2 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_2 <= trans_io_next_reg_2; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_3 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_3 <= trans_io_next_reg_3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_4 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_4 <= trans_io_next_reg_4; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_5 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_5 <= trans_io_next_reg_5; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_6 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_6 <= trans_io_next_reg_6; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_7 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_7 <= trans_io_next_reg_7; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_8 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_8 <= trans_io_next_reg_8; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_9 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_9 <= trans_io_next_reg_9; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_10 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_10 <= trans_io_next_reg_10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_11 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_11 <= trans_io_next_reg_11; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_12 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_12 <= trans_io_next_reg_12; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_13 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_13 <= trans_io_next_reg_13; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_14 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_14 <= trans_io_next_reg_14; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_15 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_15 <= trans_io_next_reg_15; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_16 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_16 <= trans_io_next_reg_16; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_17 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_17 <= trans_io_next_reg_17; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_18 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_18 <= trans_io_next_reg_18; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_19 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_19 <= trans_io_next_reg_19; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_20 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_20 <= trans_io_next_reg_20; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_21 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_21 <= trans_io_next_reg_21; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_22 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_22 <= trans_io_next_reg_22; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_23 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_23 <= trans_io_next_reg_23; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_24 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_24 <= trans_io_next_reg_24; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_25 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_25 <= trans_io_next_reg_25; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_26 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_26 <= trans_io_next_reg_26; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_27 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_27 <= trans_io_next_reg_27; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_28 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_28 <= trans_io_next_reg_28; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_29 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_29 <= trans_io_next_reg_29; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_30 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_30 <= trans_io_next_reg_30; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_reg_31 <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_reg_31 <= trans_io_next_reg_31; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_pc <= 64'h8000; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_pc <= trans_io_next_pc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_misa <= 64'h8000000000101105; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_misa <= trans_io_next_csr_misa; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mvendorid <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mvendorid <= trans_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_marchid <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_marchid <= trans_io_next_csr_marchid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mimpid <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mimpid <= trans_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mhartid <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mhartid <= trans_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mstatus <= 64'h1800; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mstatus <= trans_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mscratch <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mscratch <= trans_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mtvec <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mtvec <= trans_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mcounteren <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mcounteren <= trans_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_medeleg <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_medeleg <= trans_io_next_csr_medeleg; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mip <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mip <= trans_io_next_csr_mip; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mie <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mie <= trans_io_next_csr_mie; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mepc <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mepc <= trans_io_next_csr_mepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mcause <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mcause <= trans_io_next_csr_mcause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_mtval <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_mtval <= trans_io_next_csr_mtval; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_scause <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_scause <= trans_io_next_csr_scause; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_stvec <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_stvec <= trans_io_next_csr_stvec; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_sepc <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_sepc <= trans_io_next_csr_sepc; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_satp <= 64'h0; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_satp <= trans_io_next_csr_satp; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_MXLEN <= 8'h40; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_MXLEN <= trans_io_next_csr_MXLEN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_csr_IALIGN <= 8'h10; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_csr_IALIGN <= trans_io_next_csr_IALIGN; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
    if (reset) begin // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
      state_internal_privilegeMode <= 2'h3; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 189:22]
    end else begin
      state_internal_privilegeMode <= trans_io_next_internal_privilegeMode; // @[src/main/scala/rvspeccore/core/RiscvCore.scala 198:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  state_reg_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  state_reg_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  state_reg_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  state_reg_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  state_reg_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  state_reg_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  state_reg_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  state_reg_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  state_reg_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  state_reg_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  state_reg_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  state_reg_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  state_reg_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  state_reg_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  state_reg_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  state_reg_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  state_reg_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  state_reg_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  state_reg_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  state_reg_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  state_reg_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  state_reg_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  state_reg_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  state_reg_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  state_reg_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  state_reg_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  state_reg_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  state_reg_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  state_reg_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  state_reg_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  state_reg_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  state_reg_31 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  state_pc = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  state_csr_misa = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  state_csr_mvendorid = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  state_csr_marchid = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  state_csr_mimpid = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  state_csr_mhartid = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  state_csr_mstatus = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  state_csr_mscratch = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  state_csr_mtvec = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  state_csr_mcounteren = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  state_csr_medeleg = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  state_csr_mip = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  state_csr_mie = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  state_csr_mepc = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  state_csr_mcause = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  state_csr_mtval = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  state_csr_scause = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  state_csr_stvec = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  state_csr_sepc = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  state_csr_satp = _RAND_51[63:0];
  _RAND_52 = {1{`RANDOM}};
  state_csr_MXLEN = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  state_csr_IALIGN = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  state_internal_privilegeMode = _RAND_54[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  input  [63:0] io_enq_bits_addr, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  input  [63:0] io_enq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  output [63:0] io_deq_bits_addr, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  output [63:0] io_deq_bits_data // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_addr [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [63:0] ram_addr_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [63:0] ram_addr_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_addr_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_addr_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_addr_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  reg [63:0] ram_data [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [63:0] ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_data_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_data_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_data_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  reg  enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 277:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 278:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 279:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 280:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 304:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 303:19]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 311:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 311:17]
  always @(posedge clock) begin
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 287:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 291:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 277:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 277:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 294:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 295:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module QueueModuleTLB(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 43:14]
  input  [63:0] io_in_bits_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 43:14]
  input  [63:0] io_in_bits_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 43:14]
  input         io_out_ready, // @[src/main/scala/rvspeccore/checker/Checker.scala 43:14]
  output [63:0] io_out_bits_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 43:14]
  output [63:0] io_out_bits_data // @[src/main/scala/rvspeccore/checker/Checker.scala 43:14]
);
  wire  queue_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire  queue_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire  queue_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire  queue_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire [63:0] queue_q_io_enq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire [63:0] queue_q_io_enq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire  queue_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire  queue_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire [63:0] queue_q_io_deq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire [63:0] queue_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  Queue queue_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
    .clock(queue_q_clock),
    .reset(queue_q_reset),
    .io_enq_ready(queue_q_io_enq_ready),
    .io_enq_valid(queue_q_io_enq_valid),
    .io_enq_bits_addr(queue_q_io_enq_bits_addr),
    .io_enq_bits_data(queue_q_io_enq_bits_data),
    .io_deq_ready(queue_q_io_deq_ready),
    .io_deq_valid(queue_q_io_deq_valid),
    .io_deq_bits_addr(queue_q_io_deq_bits_addr),
    .io_deq_bits_data(queue_q_io_deq_bits_data)
  );
  assign io_out_bits_addr = queue_q_io_deq_bits_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 49:10]
  assign io_out_bits_data = queue_q_io_deq_bits_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 49:10]
  assign queue_q_clock = clock;
  assign queue_q_reset = reset;
  assign queue_q_io_enq_valid = io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 378:22]
  assign queue_q_io_enq_bits_addr = io_in_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 379:21]
  assign queue_q_io_enq_bits_data = io_in_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 379:21]
  assign queue_q_io_deq_ready = io_out_ready; // @[src/main/scala/rvspeccore/checker/Checker.scala 49:10]
endmodule
module Queue_3(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  input  [63:0] io_enq_bits_addr, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  input  [63:0] io_enq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  input  [6:0]  io_enq_bits_memWidth, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  output [63:0] io_deq_bits_addr, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  output [63:0] io_deq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
  output [6:0]  io_deq_bits_memWidth // @[src/main/scala/chisel3/util/Decoupled.scala 273:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_addr [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [63:0] ram_addr_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [63:0] ram_addr_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_addr_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_addr_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_addr_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  reg [63:0] ram_data [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [63:0] ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_data_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_data_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_data_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  reg [6:0] ram_memWidth [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_memWidth_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_memWidth_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [6:0] ram_memWidth_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire [6:0] ram_memWidth_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_memWidth_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_memWidth_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  wire  ram_memWidth_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  reg  enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 277:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 278:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 279:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 280:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_memWidth_io_deq_bits_MPORT_en = 1'h1;
  assign ram_memWidth_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_memWidth_io_deq_bits_MPORT_data = ram_memWidth[ram_memWidth_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
  assign ram_memWidth_MPORT_data = io_enq_bits_memWidth;
  assign ram_memWidth_MPORT_addr = enq_ptr_value;
  assign ram_memWidth_MPORT_mask = 1'h1;
  assign ram_memWidth_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 304:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 303:19]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 311:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 311:17]
  assign io_deq_bits_memWidth = ram_memWidth_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 311:17]
  always @(posedge clock) begin
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
    end
    if (ram_memWidth_MPORT_en & ram_memWidth_MPORT_mask) begin
      ram_memWidth[ram_memWidth_MPORT_addr] <= ram_memWidth_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 274:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 287:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 291:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 277:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 277:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 294:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 295:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_memWidth[initvar] = _RAND_2[6:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enq_ptr_value = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  deq_ptr_value = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module QueueModule(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 34:14]
  input  [63:0] io_in_bits_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 34:14]
  input  [63:0] io_in_bits_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 34:14]
  input  [6:0]  io_in_bits_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 34:14]
  input         io_out_ready, // @[src/main/scala/rvspeccore/checker/Checker.scala 34:14]
  output [63:0] io_out_bits_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 34:14]
  output [63:0] io_out_bits_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 34:14]
  output [6:0]  io_out_bits_memWidth // @[src/main/scala/rvspeccore/checker/Checker.scala 34:14]
);
  wire  queue_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire  queue_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire  queue_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire  queue_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire [63:0] queue_q_io_enq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire [63:0] queue_q_io_enq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire [6:0] queue_q_io_enq_bits_memWidth; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire  queue_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire  queue_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire [63:0] queue_q_io_deq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire [63:0] queue_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  wire [6:0] queue_q_io_deq_bits_memWidth; // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
  Queue_3 queue_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 376:21]
    .clock(queue_q_clock),
    .reset(queue_q_reset),
    .io_enq_ready(queue_q_io_enq_ready),
    .io_enq_valid(queue_q_io_enq_valid),
    .io_enq_bits_addr(queue_q_io_enq_bits_addr),
    .io_enq_bits_data(queue_q_io_enq_bits_data),
    .io_enq_bits_memWidth(queue_q_io_enq_bits_memWidth),
    .io_deq_ready(queue_q_io_deq_ready),
    .io_deq_valid(queue_q_io_deq_valid),
    .io_deq_bits_addr(queue_q_io_deq_bits_addr),
    .io_deq_bits_data(queue_q_io_deq_bits_data),
    .io_deq_bits_memWidth(queue_q_io_deq_bits_memWidth)
  );
  assign io_out_bits_addr = queue_q_io_deq_bits_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 40:10]
  assign io_out_bits_data = queue_q_io_deq_bits_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 40:10]
  assign io_out_bits_memWidth = queue_q_io_deq_bits_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 40:10]
  assign queue_q_clock = clock;
  assign queue_q_reset = reset;
  assign queue_q_io_enq_valid = io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 378:22]
  assign queue_q_io_enq_bits_addr = io_in_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 379:21]
  assign queue_q_io_enq_bits_data = io_in_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 379:21]
  assign queue_q_io_enq_bits_memWidth = io_in_bits_memWidth; // @[src/main/scala/chisel3/util/Decoupled.scala 379:21]
  assign queue_q_io_deq_ready = io_out_ready; // @[src/main/scala/rvspeccore/checker/Checker.scala 40:10]
endmodule
module CheckerWithResult(
  input         clock,
  input         reset,
  input         io_instCommit_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [31:0] io_instCommit_inst, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_instCommit_pc, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_0, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_1, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_2, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_3, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_4, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_5, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_6, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_7, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_8, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_9, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_10, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_11, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_12, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_13, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_14, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_15, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_16, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_17, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_18, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_19, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_20, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_21, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_22, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_23, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_24, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_25, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_26, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_27, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_28, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_29, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_30, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_reg_31, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_misa, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mvendorid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_marchid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mimpid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mhartid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mstatus, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mscratch, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mtvec, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mcounteren, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mip, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mie, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mepc, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mcause, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_result_csr_mtval, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input         io_event_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_event_intrNO, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_event_cause, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_event_exceptionPC, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_event_exceptionInst, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input         io_mem_read_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_mem_read_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [6:0]  io_mem_read_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_mem_read_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input         io_mem_write_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_mem_write_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [6:0]  io_mem_write_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_mem_write_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input         io_dtlbmem_read_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_dtlbmem_read_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [63:0] io_dtlbmem_read_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
  input  [1:0]  io_dtlbmem_read_level // @[src/main/scala/rvspeccore/checker/Checker.scala 63:16]
);
  wire  specCore_clock; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire  specCore_reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [31:0] specCore_io_inst; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire  specCore_io_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire  specCore_io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_mem_read_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [6:0] specCore_io_mem_read_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_mem_read_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire  specCore_io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_mem_write_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [6:0] specCore_io_mem_write_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_mem_write_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire  specCore_io_tlb_Anotherread_0_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_tlb_Anotherread_0_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_tlb_Anotherread_0_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire  specCore_io_tlb_Anotherread_1_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_tlb_Anotherread_1_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_tlb_Anotherread_1_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire  specCore_io_tlb_Anotherread_2_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_tlb_Anotherread_2_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_tlb_Anotherread_2_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_now_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_0; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_1; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_3; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_4; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_6; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_7; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_8; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_9; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_10; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_11; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_12; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_13; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_14; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_15; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_16; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_17; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_18; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_19; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_20; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_21; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_22; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_23; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_24; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_25; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_26; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_27; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_28; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_29; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_30; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_reg_31; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_misa; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mvendorid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_marchid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mimpid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mhartid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mstatus; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mtvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mcounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mip; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mie; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mcause; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_next_csr_mtval; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire  specCore_io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_event_cause; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_event_exceptionPC; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire [63:0] specCore_io_event_exceptionInst; // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
  wire  TLBLoadQueue_0_clock; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire  TLBLoadQueue_0_reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire  TLBLoadQueue_0_io_in_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire [63:0] TLBLoadQueue_0_io_in_bits_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire [63:0] TLBLoadQueue_0_io_in_bits_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire  TLBLoadQueue_0_io_out_ready; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire [63:0] TLBLoadQueue_0_io_out_bits_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire [63:0] TLBLoadQueue_0_io_out_bits_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire  TLBLoadQueue_1_clock; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire  TLBLoadQueue_1_reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire  TLBLoadQueue_1_io_in_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire [63:0] TLBLoadQueue_1_io_in_bits_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire [63:0] TLBLoadQueue_1_io_in_bits_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire  TLBLoadQueue_1_io_out_ready; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire [63:0] TLBLoadQueue_1_io_out_bits_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire [63:0] TLBLoadQueue_1_io_out_bits_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire  TLBLoadQueue_2_clock; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire  TLBLoadQueue_2_reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire  TLBLoadQueue_2_io_in_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire [63:0] TLBLoadQueue_2_io_in_bits_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire [63:0] TLBLoadQueue_2_io_in_bits_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire  TLBLoadQueue_2_io_out_ready; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire [63:0] TLBLoadQueue_2_io_out_bits_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire [63:0] TLBLoadQueue_2_io_out_bits_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
  wire  LoadQueue_clock; // @[src/main/scala/rvspeccore/checker/Checker.scala 147:30]
  wire  LoadQueue_reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 147:30]
  wire  LoadQueue_io_in_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 147:30]
  wire [63:0] LoadQueue_io_in_bits_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 147:30]
  wire [63:0] LoadQueue_io_in_bits_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 147:30]
  wire [6:0] LoadQueue_io_in_bits_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 147:30]
  wire  LoadQueue_io_out_ready; // @[src/main/scala/rvspeccore/checker/Checker.scala 147:30]
  wire [63:0] LoadQueue_io_out_bits_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 147:30]
  wire [63:0] LoadQueue_io_out_bits_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 147:30]
  wire [6:0] LoadQueue_io_out_bits_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 147:30]
  wire  StoreQueue_clock; // @[src/main/scala/rvspeccore/checker/Checker.scala 148:30]
  wire  StoreQueue_reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 148:30]
  wire  StoreQueue_io_in_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 148:30]
  wire [63:0] StoreQueue_io_in_bits_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 148:30]
  wire [63:0] StoreQueue_io_in_bits_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 148:30]
  wire [6:0] StoreQueue_io_in_bits_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 148:30]
  wire  StoreQueue_io_out_ready; // @[src/main/scala/rvspeccore/checker/Checker.scala 148:30]
  wire [63:0] StoreQueue_io_out_bits_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 148:30]
  wire [63:0] StoreQueue_io_out_bits_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 148:30]
  wire [6:0] StoreQueue_io_out_bits_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 148:30]
  wire  _T = io_dtlbmem_read_level == 2'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 127:42]
  wire [63:0] _GEN_1 = io_dtlbmem_read_level == 2'h0 ? io_dtlbmem_read_addr : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 122:38 127:51 129:46]
  wire [63:0] _GEN_2 = io_dtlbmem_read_level == 2'h0 ? io_dtlbmem_read_data : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 122:38 127:51 130:46]
  wire  _T_1 = io_dtlbmem_read_level == 2'h1; // @[src/main/scala/rvspeccore/checker/Checker.scala 127:42]
  wire [63:0] _GEN_5 = io_dtlbmem_read_level == 2'h1 ? io_dtlbmem_read_addr : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 122:38 127:51 129:46]
  wire [63:0] _GEN_6 = io_dtlbmem_read_level == 2'h1 ? io_dtlbmem_read_data : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 122:38 127:51 130:46]
  wire  _T_2 = io_dtlbmem_read_level == 2'h2; // @[src/main/scala/rvspeccore/checker/Checker.scala 127:42]
  wire [63:0] _GEN_9 = io_dtlbmem_read_level == 2'h2 ? io_dtlbmem_read_addr : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 122:38 127:51 129:46]
  wire [63:0] _GEN_10 = io_dtlbmem_read_level == 2'h2 ? io_dtlbmem_read_data : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 122:38 127:51 130:46]
  wire  _T_5 = ~reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 144:17]
  wire  _T_223 = io_event_valid | specCore_io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 212:33]
  wire  _T_224 = io_event_valid == specCore_io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 214:32]
  wire  _GEN_50 = specCore_io_mem_read_valid & _T_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 164:15]
  wire  _GEN_56 = specCore_io_mem_write_valid & _T_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 185:15]
  wire  _GEN_65 = io_instCommit_valid & _T_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 198:11]
  wire  _GEN_206 = _T_223 & _T_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 213:11]
  RiscvCore specCore ( // @[src/main/scala/rvspeccore/checker/Checker.scala 87:24]
    .clock(specCore_clock),
    .reset(specCore_reset),
    .io_inst(specCore_io_inst),
    .io_valid(specCore_io_valid),
    .io_mem_read_valid(specCore_io_mem_read_valid),
    .io_mem_read_addr(specCore_io_mem_read_addr),
    .io_mem_read_memWidth(specCore_io_mem_read_memWidth),
    .io_mem_read_data(specCore_io_mem_read_data),
    .io_mem_write_valid(specCore_io_mem_write_valid),
    .io_mem_write_addr(specCore_io_mem_write_addr),
    .io_mem_write_memWidth(specCore_io_mem_write_memWidth),
    .io_mem_write_data(specCore_io_mem_write_data),
    .io_tlb_Anotherread_0_valid(specCore_io_tlb_Anotherread_0_valid),
    .io_tlb_Anotherread_0_addr(specCore_io_tlb_Anotherread_0_addr),
    .io_tlb_Anotherread_0_data(specCore_io_tlb_Anotherread_0_data),
    .io_tlb_Anotherread_1_valid(specCore_io_tlb_Anotherread_1_valid),
    .io_tlb_Anotherread_1_addr(specCore_io_tlb_Anotherread_1_addr),
    .io_tlb_Anotherread_1_data(specCore_io_tlb_Anotherread_1_data),
    .io_tlb_Anotherread_2_valid(specCore_io_tlb_Anotherread_2_valid),
    .io_tlb_Anotherread_2_addr(specCore_io_tlb_Anotherread_2_addr),
    .io_tlb_Anotherread_2_data(specCore_io_tlb_Anotherread_2_data),
    .io_now_pc(specCore_io_now_pc),
    .io_next_reg_0(specCore_io_next_reg_0),
    .io_next_reg_1(specCore_io_next_reg_1),
    .io_next_reg_2(specCore_io_next_reg_2),
    .io_next_reg_3(specCore_io_next_reg_3),
    .io_next_reg_4(specCore_io_next_reg_4),
    .io_next_reg_5(specCore_io_next_reg_5),
    .io_next_reg_6(specCore_io_next_reg_6),
    .io_next_reg_7(specCore_io_next_reg_7),
    .io_next_reg_8(specCore_io_next_reg_8),
    .io_next_reg_9(specCore_io_next_reg_9),
    .io_next_reg_10(specCore_io_next_reg_10),
    .io_next_reg_11(specCore_io_next_reg_11),
    .io_next_reg_12(specCore_io_next_reg_12),
    .io_next_reg_13(specCore_io_next_reg_13),
    .io_next_reg_14(specCore_io_next_reg_14),
    .io_next_reg_15(specCore_io_next_reg_15),
    .io_next_reg_16(specCore_io_next_reg_16),
    .io_next_reg_17(specCore_io_next_reg_17),
    .io_next_reg_18(specCore_io_next_reg_18),
    .io_next_reg_19(specCore_io_next_reg_19),
    .io_next_reg_20(specCore_io_next_reg_20),
    .io_next_reg_21(specCore_io_next_reg_21),
    .io_next_reg_22(specCore_io_next_reg_22),
    .io_next_reg_23(specCore_io_next_reg_23),
    .io_next_reg_24(specCore_io_next_reg_24),
    .io_next_reg_25(specCore_io_next_reg_25),
    .io_next_reg_26(specCore_io_next_reg_26),
    .io_next_reg_27(specCore_io_next_reg_27),
    .io_next_reg_28(specCore_io_next_reg_28),
    .io_next_reg_29(specCore_io_next_reg_29),
    .io_next_reg_30(specCore_io_next_reg_30),
    .io_next_reg_31(specCore_io_next_reg_31),
    .io_next_csr_misa(specCore_io_next_csr_misa),
    .io_next_csr_mvendorid(specCore_io_next_csr_mvendorid),
    .io_next_csr_marchid(specCore_io_next_csr_marchid),
    .io_next_csr_mimpid(specCore_io_next_csr_mimpid),
    .io_next_csr_mhartid(specCore_io_next_csr_mhartid),
    .io_next_csr_mstatus(specCore_io_next_csr_mstatus),
    .io_next_csr_mscratch(specCore_io_next_csr_mscratch),
    .io_next_csr_mtvec(specCore_io_next_csr_mtvec),
    .io_next_csr_mcounteren(specCore_io_next_csr_mcounteren),
    .io_next_csr_mip(specCore_io_next_csr_mip),
    .io_next_csr_mie(specCore_io_next_csr_mie),
    .io_next_csr_mepc(specCore_io_next_csr_mepc),
    .io_next_csr_mcause(specCore_io_next_csr_mcause),
    .io_next_csr_mtval(specCore_io_next_csr_mtval),
    .io_event_valid(specCore_io_event_valid),
    .io_event_cause(specCore_io_event_cause),
    .io_event_exceptionPC(specCore_io_event_exceptionPC),
    .io_event_exceptionInst(specCore_io_event_exceptionInst)
  );
  QueueModuleTLB TLBLoadQueue_0 ( // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
    .clock(TLBLoadQueue_0_clock),
    .reset(TLBLoadQueue_0_reset),
    .io_in_valid(TLBLoadQueue_0_io_in_valid),
    .io_in_bits_addr(TLBLoadQueue_0_io_in_bits_addr),
    .io_in_bits_data(TLBLoadQueue_0_io_in_bits_data),
    .io_out_ready(TLBLoadQueue_0_io_out_ready),
    .io_out_bits_addr(TLBLoadQueue_0_io_out_bits_addr),
    .io_out_bits_data(TLBLoadQueue_0_io_out_bits_data)
  );
  QueueModuleTLB TLBLoadQueue_1 ( // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
    .clock(TLBLoadQueue_1_clock),
    .reset(TLBLoadQueue_1_reset),
    .io_in_valid(TLBLoadQueue_1_io_in_valid),
    .io_in_bits_addr(TLBLoadQueue_1_io_in_bits_addr),
    .io_in_bits_data(TLBLoadQueue_1_io_in_bits_data),
    .io_out_ready(TLBLoadQueue_1_io_out_ready),
    .io_out_bits_addr(TLBLoadQueue_1_io_out_bits_addr),
    .io_out_bits_data(TLBLoadQueue_1_io_out_bits_data)
  );
  QueueModuleTLB TLBLoadQueue_2 ( // @[src/main/scala/rvspeccore/checker/Checker.scala 117:44]
    .clock(TLBLoadQueue_2_clock),
    .reset(TLBLoadQueue_2_reset),
    .io_in_valid(TLBLoadQueue_2_io_in_valid),
    .io_in_bits_addr(TLBLoadQueue_2_io_in_bits_addr),
    .io_in_bits_data(TLBLoadQueue_2_io_in_bits_data),
    .io_out_ready(TLBLoadQueue_2_io_out_ready),
    .io_out_bits_addr(TLBLoadQueue_2_io_out_bits_addr),
    .io_out_bits_data(TLBLoadQueue_2_io_out_bits_data)
  );
  QueueModule LoadQueue ( // @[src/main/scala/rvspeccore/checker/Checker.scala 147:30]
    .clock(LoadQueue_clock),
    .reset(LoadQueue_reset),
    .io_in_valid(LoadQueue_io_in_valid),
    .io_in_bits_addr(LoadQueue_io_in_bits_addr),
    .io_in_bits_data(LoadQueue_io_in_bits_data),
    .io_in_bits_memWidth(LoadQueue_io_in_bits_memWidth),
    .io_out_ready(LoadQueue_io_out_ready),
    .io_out_bits_addr(LoadQueue_io_out_bits_addr),
    .io_out_bits_data(LoadQueue_io_out_bits_data),
    .io_out_bits_memWidth(LoadQueue_io_out_bits_memWidth)
  );
  QueueModule StoreQueue ( // @[src/main/scala/rvspeccore/checker/Checker.scala 148:30]
    .clock(StoreQueue_clock),
    .reset(StoreQueue_reset),
    .io_in_valid(StoreQueue_io_in_valid),
    .io_in_bits_addr(StoreQueue_io_in_bits_addr),
    .io_in_bits_data(StoreQueue_io_in_bits_data),
    .io_in_bits_memWidth(StoreQueue_io_in_bits_memWidth),
    .io_out_ready(StoreQueue_io_out_ready),
    .io_out_bits_addr(StoreQueue_io_out_bits_addr),
    .io_out_bits_data(StoreQueue_io_out_bits_data),
    .io_out_bits_memWidth(StoreQueue_io_out_bits_memWidth)
  );
  assign specCore_clock = clock;
  assign specCore_reset = reset;
  assign specCore_io_inst = io_instCommit_inst; // @[src/main/scala/rvspeccore/checker/Checker.scala 89:21]
  assign specCore_io_valid = io_instCommit_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 88:21]
  assign specCore_io_mem_read_data = specCore_io_mem_read_valid ? LoadQueue_io_out_bits_data : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 160:50 163:35 168:35]
  assign specCore_io_tlb_Anotherread_0_data = TLBLoadQueue_2_io_out_bits_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 136:56 139:51]
  assign specCore_io_tlb_Anotherread_1_data = TLBLoadQueue_1_io_out_bits_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 136:56 139:51]
  assign specCore_io_tlb_Anotherread_2_data = TLBLoadQueue_0_io_out_bits_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 136:56 139:51]
  assign TLBLoadQueue_0_clock = clock;
  assign TLBLoadQueue_0_reset = reset;
  assign TLBLoadQueue_0_io_in_valid = io_dtlbmem_read_valid & _T; // @[src/main/scala/rvspeccore/checker/Checker.scala 121:38 124:39]
  assign TLBLoadQueue_0_io_in_bits_addr = io_dtlbmem_read_valid ? _GEN_1 : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 122:38 124:39]
  assign TLBLoadQueue_0_io_in_bits_data = io_dtlbmem_read_valid ? _GEN_2 : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 122:38 124:39]
  assign TLBLoadQueue_0_io_out_ready = specCore_io_tlb_Anotherread_2_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 120:38 136:56 137:44]
  assign TLBLoadQueue_1_clock = clock;
  assign TLBLoadQueue_1_reset = reset;
  assign TLBLoadQueue_1_io_in_valid = io_dtlbmem_read_valid & _T_1; // @[src/main/scala/rvspeccore/checker/Checker.scala 121:38 124:39]
  assign TLBLoadQueue_1_io_in_bits_addr = io_dtlbmem_read_valid ? _GEN_5 : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 122:38 124:39]
  assign TLBLoadQueue_1_io_in_bits_data = io_dtlbmem_read_valid ? _GEN_6 : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 122:38 124:39]
  assign TLBLoadQueue_1_io_out_ready = specCore_io_tlb_Anotherread_1_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 120:38 136:56 137:44]
  assign TLBLoadQueue_2_clock = clock;
  assign TLBLoadQueue_2_reset = reset;
  assign TLBLoadQueue_2_io_in_valid = io_dtlbmem_read_valid & _T_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 121:38 124:39]
  assign TLBLoadQueue_2_io_in_bits_addr = io_dtlbmem_read_valid ? _GEN_9 : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 122:38 124:39]
  assign TLBLoadQueue_2_io_in_bits_data = io_dtlbmem_read_valid ? _GEN_10 : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 122:38 124:39]
  assign TLBLoadQueue_2_io_out_ready = specCore_io_tlb_Anotherread_0_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 120:38 136:56 137:44]
  assign LoadQueue_clock = clock;
  assign LoadQueue_reset = reset;
  assign LoadQueue_io_in_valid = io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 150:35 151:39 157:31]
  assign LoadQueue_io_in_bits_addr = io_mem_read_valid ? io_mem_read_addr : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 150:35 152:39 158:31]
  assign LoadQueue_io_in_bits_data = io_mem_read_valid ? io_mem_read_data : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 150:35 153:39 158:31]
  assign LoadQueue_io_in_bits_memWidth = io_mem_read_valid ? io_mem_read_memWidth : 7'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 150:35 154:39 158:31]
  assign LoadQueue_io_out_ready = specCore_io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 160:50 161:32 167:35]
  assign StoreQueue_clock = clock;
  assign StoreQueue_reset = reset;
  assign StoreQueue_io_in_valid = io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 172:36 173:40 179:32]
  assign StoreQueue_io_in_bits_addr = io_mem_write_valid ? io_mem_write_addr : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 172:36 174:40 180:32]
  assign StoreQueue_io_in_bits_data = io_mem_write_valid ? io_mem_write_data : 64'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 172:36 175:40 180:32]
  assign StoreQueue_io_in_bits_memWidth = io_mem_write_valid ? io_mem_write_memWidth : 7'h0; // @[src/main/scala/rvspeccore/checker/Checker.scala 172:36 176:40 180:32]
  assign StoreQueue_io_out_ready = specCore_io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 182:51 183:33 189:33]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (specCore_io_tlb_Anotherread_0_valid & ~reset & ~(TLBLoadQueue_2_io_out_bits_addr ==
          specCore_io_tlb_Anotherread_0_addr)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:144 assert(regDelay(TLBLoadQueue(2 - i).io.out.bits.addr) === regDelay(specCore.io.tlb.get.Anotherread(i).addr))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 144:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (specCore_io_tlb_Anotherread_0_valid & ~reset & ~(TLBLoadQueue_2_io_out_bits_addr ==
          specCore_io_tlb_Anotherread_0_addr)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 144:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (specCore_io_tlb_Anotherread_1_valid & ~reset & ~(TLBLoadQueue_1_io_out_bits_addr ==
          specCore_io_tlb_Anotherread_1_addr)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:144 assert(regDelay(TLBLoadQueue(2 - i).io.out.bits.addr) === regDelay(specCore.io.tlb.get.Anotherread(i).addr))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 144:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (specCore_io_tlb_Anotherread_1_valid & ~reset & ~(TLBLoadQueue_1_io_out_bits_addr ==
          specCore_io_tlb_Anotherread_1_addr)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 144:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (specCore_io_tlb_Anotherread_2_valid & ~reset & ~(TLBLoadQueue_0_io_out_bits_addr ==
          specCore_io_tlb_Anotherread_2_addr)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:144 assert(regDelay(TLBLoadQueue(2 - i).io.out.bits.addr) === regDelay(specCore.io.tlb.get.Anotherread(i).addr))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 144:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (specCore_io_tlb_Anotherread_2_valid & ~reset & ~(TLBLoadQueue_0_io_out_bits_addr ==
          specCore_io_tlb_Anotherread_2_addr)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 144:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (specCore_io_mem_read_valid & _T_5 & ~(LoadQueue_io_out_bits_addr == specCore_io_mem_read_addr)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:164 assert(regDelay(LoadQueue.io.out.bits.addr) === regDelay(specCore.io.mem.read.addr))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 164:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (specCore_io_mem_read_valid & _T_5 & ~(LoadQueue_io_out_bits_addr == specCore_io_mem_read_addr)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 164:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_50 & ~(LoadQueue_io_out_bits_memWidth == specCore_io_mem_read_memWidth)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:165 assert(regDelay(LoadQueue.io.out.bits.memWidth) === regDelay(specCore.io.mem.read.memWidth))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 165:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_50 & ~(LoadQueue_io_out_bits_memWidth == specCore_io_mem_read_memWidth)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 165:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (specCore_io_mem_write_valid & _T_5 & ~(StoreQueue_io_out_bits_addr == specCore_io_mem_write_addr)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:185 assert(regDelay(StoreQueue.io.out.bits.addr) === regDelay(specCore.io.mem.write.addr))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 185:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (specCore_io_mem_write_valid & _T_5 & ~(StoreQueue_io_out_bits_addr == specCore_io_mem_write_addr)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 185:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & ~(StoreQueue_io_out_bits_data == specCore_io_mem_write_data)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:186 assert(regDelay(StoreQueue.io.out.bits.data) === regDelay(specCore.io.mem.write.data))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 186:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_56 & ~(StoreQueue_io_out_bits_data == specCore_io_mem_write_data)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 186:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & ~(StoreQueue_io_out_bits_memWidth == specCore_io_mem_write_memWidth)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:187 assert(regDelay(StoreQueue.io.out.bits.memWidth) === regDelay(specCore.io.mem.write.memWidth))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 187:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_56 & ~(StoreQueue_io_out_bits_memWidth == specCore_io_mem_write_memWidth)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 187:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_instCommit_valid & _T_5 & ~(io_instCommit_pc == specCore_io_now_pc)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:198 assert(regDelay(io.instCommit.pc) === regDelay(specCore.io.now.pc))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 198:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_instCommit_valid & _T_5 & ~(io_instCommit_pc == specCore_io_now_pc)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 198:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_misa == specCore_io_next_csr_misa)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_misa == specCore_io_next_csr_misa)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mvendorid == specCore_io_next_csr_mvendorid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mvendorid == specCore_io_next_csr_mvendorid)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_marchid == specCore_io_next_csr_marchid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_marchid == specCore_io_next_csr_marchid)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mimpid == specCore_io_next_csr_mimpid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mimpid == specCore_io_next_csr_mimpid)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mhartid == specCore_io_next_csr_mhartid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mhartid == specCore_io_next_csr_mhartid)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mstatus == specCore_io_next_csr_mstatus)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mstatus == specCore_io_next_csr_mstatus)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mscratch == specCore_io_next_csr_mscratch)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mscratch == specCore_io_next_csr_mscratch)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mtvec == specCore_io_next_csr_mtvec)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mtvec == specCore_io_next_csr_mtvec)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mcounteren == specCore_io_next_csr_mcounteren)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mcounteren == specCore_io_next_csr_mcounteren)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mip == specCore_io_next_csr_mip)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mip == specCore_io_next_csr_mip)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mie == specCore_io_next_csr_mie)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mie == specCore_io_next_csr_mie)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mepc == specCore_io_next_csr_mepc)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mepc == specCore_io_next_csr_mepc)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mcause == specCore_io_next_csr_mcause)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mcause == specCore_io_next_csr_mcause)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mtval == specCore_io_next_csr_mtval)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:203 assert(regDelay(result.signal) === regDelay(next.signal))\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_csr_mtval == specCore_io_next_csr_mtval)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 203:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_0 == specCore_io_next_reg_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_0 == specCore_io_next_reg_0)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_1 == specCore_io_next_reg_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_1 == specCore_io_next_reg_1)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_2 == specCore_io_next_reg_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_2 == specCore_io_next_reg_2)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_3 == specCore_io_next_reg_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_3 == specCore_io_next_reg_3)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_4 == specCore_io_next_reg_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_4 == specCore_io_next_reg_4)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_5 == specCore_io_next_reg_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_5 == specCore_io_next_reg_5)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_6 == specCore_io_next_reg_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_6 == specCore_io_next_reg_6)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_7 == specCore_io_next_reg_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_7 == specCore_io_next_reg_7)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_8 == specCore_io_next_reg_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_8 == specCore_io_next_reg_8)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_9 == specCore_io_next_reg_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_9 == specCore_io_next_reg_9)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_10 == specCore_io_next_reg_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_10 == specCore_io_next_reg_10)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_11 == specCore_io_next_reg_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_11 == specCore_io_next_reg_11)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_12 == specCore_io_next_reg_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_12 == specCore_io_next_reg_12)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_13 == specCore_io_next_reg_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_13 == specCore_io_next_reg_13)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_14 == specCore_io_next_reg_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_14 == specCore_io_next_reg_14)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_15 == specCore_io_next_reg_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_15 == specCore_io_next_reg_15)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_16 == specCore_io_next_reg_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_16 == specCore_io_next_reg_16)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_17 == specCore_io_next_reg_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_17 == specCore_io_next_reg_17)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_18 == specCore_io_next_reg_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_18 == specCore_io_next_reg_18)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_19 == specCore_io_next_reg_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_19 == specCore_io_next_reg_19)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_20 == specCore_io_next_reg_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_20 == specCore_io_next_reg_20)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_21 == specCore_io_next_reg_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_21 == specCore_io_next_reg_21)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_22 == specCore_io_next_reg_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_22 == specCore_io_next_reg_22)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_23 == specCore_io_next_reg_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_23 == specCore_io_next_reg_23)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_24 == specCore_io_next_reg_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_24 == specCore_io_next_reg_24)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_25 == specCore_io_next_reg_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_25 == specCore_io_next_reg_25)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_26 == specCore_io_next_reg_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_26 == specCore_io_next_reg_26)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_27 == specCore_io_next_reg_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_27 == specCore_io_next_reg_27)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_28 == specCore_io_next_reg_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_28 == specCore_io_next_reg_28)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_29 == specCore_io_next_reg_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_29 == specCore_io_next_reg_29)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_30 == specCore_io_next_reg_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_30 == specCore_io_next_reg_30)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_31 == specCore_io_next_reg_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:208 assert(regDelay(io.result.reg(i.U)) === regDelay(specCore.io.next.reg(i.U)))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & ~(io_result_reg_31 == specCore_io_next_reg_31)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 208:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_223 & _T_5 & ~_T_224) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Checker.scala:213 assert(\n"); // @[src/main/scala/rvspeccore/checker/Checker.scala 213:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_223 & _T_5 & ~_T_224) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 213:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_206 & ~(io_event_intrNO == 64'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:216 assert(regDelay(io.event.intrNO) === regDelay(specCore.io.event.intrNO))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 216:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_206 & ~(io_event_intrNO == 64'h0)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 216:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_206 & ~(io_event_cause == specCore_io_event_cause)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:217 assert(regDelay(io.event.cause) === regDelay(specCore.io.event.cause))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 217:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_206 & ~(io_event_cause == specCore_io_event_cause)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 217:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_206 & ~(io_event_exceptionPC == specCore_io_event_exceptionPC)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:218 assert(regDelay(io.event.exceptionPC) === regDelay(specCore.io.event.exceptionPC))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 218:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_206 & ~(io_event_exceptionPC == specCore_io_event_exceptionPC)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 218:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_206 & ~(io_event_exceptionInst == specCore_io_event_exceptionInst)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Checker.scala:219 assert(regDelay(io.event.exceptionInst) === regDelay(specCore.io.event.exceptionInst))\n"
            ); // @[src/main/scala/rvspeccore/checker/Checker.scala 219:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_206 & ~(io_event_exceptionInst == specCore_io_event_exceptionInst)) begin
          $fatal; // @[src/main/scala/rvspeccore/checker/Checker.scala 219:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CheckerWrapper(
  input         clock,
  input         reset,
  input         io_instCommit_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [31:0] io_instCommit_inst, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_instCommit_pc, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_0, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_1, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_2, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_3, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_4, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_5, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_6, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_7, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_8, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_9, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_10, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_11, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_12, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_13, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_14, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_15, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_16, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_17, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_18, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_19, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_20, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_21, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_22, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_23, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_24, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_25, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_26, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_27, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_28, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_29, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_30, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_reg_31, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_pc, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_misa, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_mvendorid, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_marchid, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_mimpid, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_mhartid, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_mstatus, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_mstatush, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_mscratch, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_mtvec, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_mcounteren, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_medeleg, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_mideleg, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_mip, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_mie, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_mepc, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_mcause, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_mtval, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_cycle, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_scounteren, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_scause, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_stvec, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_sepc, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_stval, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_sscratch, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_satp, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_pmpcfg0, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_pmpcfg1, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_pmpcfg2, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_pmpcfg3, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_pmpaddr0, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_pmpaddr1, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_pmpaddr2, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_result_csr_pmpaddr3, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [7:0]  io_result_csr_MXLEN, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [7:0]  io_result_csr_IALIGN, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [7:0]  io_result_csr_ILEN, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [1:0]  io_result_internal_privilegeMode, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input         io_event_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_event_intrNO, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_event_cause, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_event_exceptionPC, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_event_exceptionInst, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input         io_mem_read_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_mem_read_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [6:0]  io_mem_read_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_mem_read_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input         io_mem_write_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_mem_write_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [6:0]  io_mem_write_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_mem_write_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input         io_dtlbmem_read_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_dtlbmem_read_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_dtlbmem_read_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [6:0]  io_dtlbmem_read_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input         io_dtlbmem_read_access, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [1:0]  io_dtlbmem_read_level, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input         io_dtlbmem_write_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_dtlbmem_write_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_dtlbmem_write_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [6:0]  io_dtlbmem_write_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input         io_dtlbmem_write_access, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [1:0]  io_dtlbmem_write_level, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input         io_itlbmem_read_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_itlbmem_read_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_itlbmem_read_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [6:0]  io_itlbmem_read_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input         io_itlbmem_read_access, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [1:0]  io_itlbmem_read_level, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input         io_itlbmem_write_valid, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_itlbmem_write_addr, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [63:0] io_itlbmem_write_data, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [6:0]  io_itlbmem_write_memWidth, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input         io_itlbmem_write_access, // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
  input  [1:0]  io_itlbmem_write_level // @[src/main/scala/rvspeccore/checker/Checker.scala 319:14]
);
  wire  checker__clock; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire  checker__reset; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire  checker__io_instCommit_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [31:0] checker__io_instCommit_inst; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_instCommit_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_0; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_1; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_3; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_4; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_6; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_7; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_8; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_9; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_10; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_11; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_12; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_13; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_14; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_15; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_16; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_17; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_18; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_19; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_20; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_21; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_22; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_23; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_24; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_25; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_26; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_27; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_28; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_29; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_30; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_reg_31; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_csr_misa; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_csr_mvendorid; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_csr_marchid; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_csr_mimpid; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_csr_mhartid; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_csr_mstatus; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_csr_mscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_csr_mtvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_csr_mcounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_csr_mip; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_csr_mie; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_csr_mepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_csr_mcause; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_result_csr_mtval; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire  checker__io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_event_intrNO; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_event_cause; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_event_exceptionPC; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_event_exceptionInst; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire  checker__io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_mem_read_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [6:0] checker__io_mem_read_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_mem_read_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire  checker__io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_mem_write_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [6:0] checker__io_mem_write_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_mem_write_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire  checker__io_dtlbmem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_dtlbmem_read_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [63:0] checker__io_dtlbmem_read_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  wire [1:0] checker__io_dtlbmem_read_level; // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
  CheckerWithResult checker_ ( // @[src/main/scala/rvspeccore/checker/Checker.scala 330:23]
    .clock(checker__clock),
    .reset(checker__reset),
    .io_instCommit_valid(checker__io_instCommit_valid),
    .io_instCommit_inst(checker__io_instCommit_inst),
    .io_instCommit_pc(checker__io_instCommit_pc),
    .io_result_reg_0(checker__io_result_reg_0),
    .io_result_reg_1(checker__io_result_reg_1),
    .io_result_reg_2(checker__io_result_reg_2),
    .io_result_reg_3(checker__io_result_reg_3),
    .io_result_reg_4(checker__io_result_reg_4),
    .io_result_reg_5(checker__io_result_reg_5),
    .io_result_reg_6(checker__io_result_reg_6),
    .io_result_reg_7(checker__io_result_reg_7),
    .io_result_reg_8(checker__io_result_reg_8),
    .io_result_reg_9(checker__io_result_reg_9),
    .io_result_reg_10(checker__io_result_reg_10),
    .io_result_reg_11(checker__io_result_reg_11),
    .io_result_reg_12(checker__io_result_reg_12),
    .io_result_reg_13(checker__io_result_reg_13),
    .io_result_reg_14(checker__io_result_reg_14),
    .io_result_reg_15(checker__io_result_reg_15),
    .io_result_reg_16(checker__io_result_reg_16),
    .io_result_reg_17(checker__io_result_reg_17),
    .io_result_reg_18(checker__io_result_reg_18),
    .io_result_reg_19(checker__io_result_reg_19),
    .io_result_reg_20(checker__io_result_reg_20),
    .io_result_reg_21(checker__io_result_reg_21),
    .io_result_reg_22(checker__io_result_reg_22),
    .io_result_reg_23(checker__io_result_reg_23),
    .io_result_reg_24(checker__io_result_reg_24),
    .io_result_reg_25(checker__io_result_reg_25),
    .io_result_reg_26(checker__io_result_reg_26),
    .io_result_reg_27(checker__io_result_reg_27),
    .io_result_reg_28(checker__io_result_reg_28),
    .io_result_reg_29(checker__io_result_reg_29),
    .io_result_reg_30(checker__io_result_reg_30),
    .io_result_reg_31(checker__io_result_reg_31),
    .io_result_csr_misa(checker__io_result_csr_misa),
    .io_result_csr_mvendorid(checker__io_result_csr_mvendorid),
    .io_result_csr_marchid(checker__io_result_csr_marchid),
    .io_result_csr_mimpid(checker__io_result_csr_mimpid),
    .io_result_csr_mhartid(checker__io_result_csr_mhartid),
    .io_result_csr_mstatus(checker__io_result_csr_mstatus),
    .io_result_csr_mscratch(checker__io_result_csr_mscratch),
    .io_result_csr_mtvec(checker__io_result_csr_mtvec),
    .io_result_csr_mcounteren(checker__io_result_csr_mcounteren),
    .io_result_csr_mip(checker__io_result_csr_mip),
    .io_result_csr_mie(checker__io_result_csr_mie),
    .io_result_csr_mepc(checker__io_result_csr_mepc),
    .io_result_csr_mcause(checker__io_result_csr_mcause),
    .io_result_csr_mtval(checker__io_result_csr_mtval),
    .io_event_valid(checker__io_event_valid),
    .io_event_intrNO(checker__io_event_intrNO),
    .io_event_cause(checker__io_event_cause),
    .io_event_exceptionPC(checker__io_event_exceptionPC),
    .io_event_exceptionInst(checker__io_event_exceptionInst),
    .io_mem_read_valid(checker__io_mem_read_valid),
    .io_mem_read_addr(checker__io_mem_read_addr),
    .io_mem_read_memWidth(checker__io_mem_read_memWidth),
    .io_mem_read_data(checker__io_mem_read_data),
    .io_mem_write_valid(checker__io_mem_write_valid),
    .io_mem_write_addr(checker__io_mem_write_addr),
    .io_mem_write_memWidth(checker__io_mem_write_memWidth),
    .io_mem_write_data(checker__io_mem_write_data),
    .io_dtlbmem_read_valid(checker__io_dtlbmem_read_valid),
    .io_dtlbmem_read_addr(checker__io_dtlbmem_read_addr),
    .io_dtlbmem_read_data(checker__io_dtlbmem_read_data),
    .io_dtlbmem_read_level(checker__io_dtlbmem_read_level)
  );
  assign checker__clock = clock;
  assign checker__reset = reset;
  assign checker__io_instCommit_valid = io_instCommit_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 333:25]
  assign checker__io_instCommit_inst = io_instCommit_inst; // @[src/main/scala/rvspeccore/checker/Checker.scala 333:25]
  assign checker__io_instCommit_pc = io_instCommit_pc; // @[src/main/scala/rvspeccore/checker/Checker.scala 333:25]
  assign checker__io_result_reg_0 = io_result_reg_0; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_1 = io_result_reg_1; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_2 = io_result_reg_2; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_3 = io_result_reg_3; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_4 = io_result_reg_4; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_5 = io_result_reg_5; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_6 = io_result_reg_6; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_7 = io_result_reg_7; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_8 = io_result_reg_8; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_9 = io_result_reg_9; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_10 = io_result_reg_10; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_11 = io_result_reg_11; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_12 = io_result_reg_12; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_13 = io_result_reg_13; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_14 = io_result_reg_14; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_15 = io_result_reg_15; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_16 = io_result_reg_16; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_17 = io_result_reg_17; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_18 = io_result_reg_18; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_19 = io_result_reg_19; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_20 = io_result_reg_20; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_21 = io_result_reg_21; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_22 = io_result_reg_22; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_23 = io_result_reg_23; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_24 = io_result_reg_24; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_25 = io_result_reg_25; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_26 = io_result_reg_26; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_27 = io_result_reg_27; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_28 = io_result_reg_28; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_29 = io_result_reg_29; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_30 = io_result_reg_30; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_reg_31 = io_result_reg_31; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_csr_misa = io_result_csr_misa; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_csr_mvendorid = io_result_csr_mvendorid; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_csr_marchid = io_result_csr_marchid; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_csr_mimpid = io_result_csr_mimpid; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_csr_mhartid = io_result_csr_mhartid; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_csr_mstatus = io_result_csr_mstatus; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_csr_mscratch = io_result_csr_mscratch; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_csr_mtvec = io_result_csr_mtvec; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_csr_mcounteren = io_result_csr_mcounteren; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_csr_mip = io_result_csr_mip; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_csr_mie = io_result_csr_mie; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_csr_mepc = io_result_csr_mepc; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_csr_mcause = io_result_csr_mcause; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_result_csr_mtval = io_result_csr_mtval; // @[src/main/scala/rvspeccore/checker/Checker.scala 334:25]
  assign checker__io_event_valid = io_event_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 335:25]
  assign checker__io_event_intrNO = io_event_intrNO; // @[src/main/scala/rvspeccore/checker/Checker.scala 335:25]
  assign checker__io_event_cause = io_event_cause; // @[src/main/scala/rvspeccore/checker/Checker.scala 335:25]
  assign checker__io_event_exceptionPC = io_event_exceptionPC; // @[src/main/scala/rvspeccore/checker/Checker.scala 335:25]
  assign checker__io_event_exceptionInst = io_event_exceptionInst; // @[src/main/scala/rvspeccore/checker/Checker.scala 335:25]
  assign checker__io_mem_read_valid = io_mem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 338:24]
  assign checker__io_mem_read_addr = io_mem_read_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 338:24]
  assign checker__io_mem_read_memWidth = io_mem_read_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 338:24]
  assign checker__io_mem_read_data = io_mem_read_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 338:24]
  assign checker__io_mem_write_valid = io_mem_write_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 338:24]
  assign checker__io_mem_write_addr = io_mem_write_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 338:24]
  assign checker__io_mem_write_memWidth = io_mem_write_memWidth; // @[src/main/scala/rvspeccore/checker/Checker.scala 338:24]
  assign checker__io_mem_write_data = io_mem_write_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 338:24]
  assign checker__io_dtlbmem_read_valid = io_dtlbmem_read_valid; // @[src/main/scala/rvspeccore/checker/Checker.scala 340:30]
  assign checker__io_dtlbmem_read_addr = io_dtlbmem_read_addr; // @[src/main/scala/rvspeccore/checker/Checker.scala 340:30]
  assign checker__io_dtlbmem_read_data = io_dtlbmem_read_data; // @[src/main/scala/rvspeccore/checker/Checker.scala 340:30]
  assign checker__io_dtlbmem_read_level = io_dtlbmem_read_level; // @[src/main/scala/rvspeccore/checker/Checker.scala 340:30]
endmodule
